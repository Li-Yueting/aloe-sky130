VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 53.600 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.965 5.085 6.435 ;
        RECT 8.315 2.965 11.785 6.435 ;
        RECT 15.015 2.965 18.485 6.435 ;
        RECT 21.715 2.965 25.185 6.435 ;
        RECT 28.415 2.965 31.885 6.435 ;
        RECT 35.115 2.965 38.585 6.435 ;
        RECT 41.815 2.965 45.285 6.435 ;
        RECT 48.515 2.965 51.985 6.435 ;
      LAYER mcon ;
        RECT 1.980 5.830 2.150 6.000 ;
        RECT 2.480 5.830 2.650 6.000 ;
        RECT 2.980 5.830 3.150 6.000 ;
        RECT 3.480 5.830 3.650 6.000 ;
        RECT 3.980 5.830 4.150 6.000 ;
        RECT 4.480 5.830 4.650 6.000 ;
        RECT 1.980 5.330 2.150 5.500 ;
        RECT 2.480 5.330 2.650 5.500 ;
        RECT 2.980 5.330 3.150 5.500 ;
        RECT 3.480 5.330 3.650 5.500 ;
        RECT 3.980 5.330 4.150 5.500 ;
        RECT 4.480 5.330 4.650 5.500 ;
        RECT 1.980 4.830 2.150 5.000 ;
        RECT 2.480 4.830 2.650 5.000 ;
        RECT 2.980 4.830 3.150 5.000 ;
        RECT 3.480 4.830 3.650 5.000 ;
        RECT 3.980 4.830 4.150 5.000 ;
        RECT 4.480 4.830 4.650 5.000 ;
        RECT 1.980 4.330 2.150 4.500 ;
        RECT 2.480 4.330 2.650 4.500 ;
        RECT 2.980 4.330 3.150 4.500 ;
        RECT 3.480 4.330 3.650 4.500 ;
        RECT 3.980 4.330 4.150 4.500 ;
        RECT 4.480 4.330 4.650 4.500 ;
        RECT 1.980 3.830 2.150 4.000 ;
        RECT 2.480 3.830 2.650 4.000 ;
        RECT 2.980 3.830 3.150 4.000 ;
        RECT 3.480 3.830 3.650 4.000 ;
        RECT 3.980 3.830 4.150 4.000 ;
        RECT 4.480 3.830 4.650 4.000 ;
        RECT 1.980 3.330 2.150 3.500 ;
        RECT 2.480 3.330 2.650 3.500 ;
        RECT 2.980 3.330 3.150 3.500 ;
        RECT 3.480 3.330 3.650 3.500 ;
        RECT 3.980 3.330 4.150 3.500 ;
        RECT 4.480 3.330 4.650 3.500 ;
        RECT 8.680 5.830 8.850 6.000 ;
        RECT 9.180 5.830 9.350 6.000 ;
        RECT 9.680 5.830 9.850 6.000 ;
        RECT 10.180 5.830 10.350 6.000 ;
        RECT 10.680 5.830 10.850 6.000 ;
        RECT 11.180 5.830 11.350 6.000 ;
        RECT 8.680 5.330 8.850 5.500 ;
        RECT 9.180 5.330 9.350 5.500 ;
        RECT 9.680 5.330 9.850 5.500 ;
        RECT 10.180 5.330 10.350 5.500 ;
        RECT 10.680 5.330 10.850 5.500 ;
        RECT 11.180 5.330 11.350 5.500 ;
        RECT 8.680 4.830 8.850 5.000 ;
        RECT 9.180 4.830 9.350 5.000 ;
        RECT 9.680 4.830 9.850 5.000 ;
        RECT 10.180 4.830 10.350 5.000 ;
        RECT 10.680 4.830 10.850 5.000 ;
        RECT 11.180 4.830 11.350 5.000 ;
        RECT 8.680 4.330 8.850 4.500 ;
        RECT 9.180 4.330 9.350 4.500 ;
        RECT 9.680 4.330 9.850 4.500 ;
        RECT 10.180 4.330 10.350 4.500 ;
        RECT 10.680 4.330 10.850 4.500 ;
        RECT 11.180 4.330 11.350 4.500 ;
        RECT 8.680 3.830 8.850 4.000 ;
        RECT 9.180 3.830 9.350 4.000 ;
        RECT 9.680 3.830 9.850 4.000 ;
        RECT 10.180 3.830 10.350 4.000 ;
        RECT 10.680 3.830 10.850 4.000 ;
        RECT 11.180 3.830 11.350 4.000 ;
        RECT 8.680 3.330 8.850 3.500 ;
        RECT 9.180 3.330 9.350 3.500 ;
        RECT 9.680 3.330 9.850 3.500 ;
        RECT 10.180 3.330 10.350 3.500 ;
        RECT 10.680 3.330 10.850 3.500 ;
        RECT 11.180 3.330 11.350 3.500 ;
        RECT 15.380 5.830 15.550 6.000 ;
        RECT 15.880 5.830 16.050 6.000 ;
        RECT 16.380 5.830 16.550 6.000 ;
        RECT 16.880 5.830 17.050 6.000 ;
        RECT 17.380 5.830 17.550 6.000 ;
        RECT 17.880 5.830 18.050 6.000 ;
        RECT 15.380 5.330 15.550 5.500 ;
        RECT 15.880 5.330 16.050 5.500 ;
        RECT 16.380 5.330 16.550 5.500 ;
        RECT 16.880 5.330 17.050 5.500 ;
        RECT 17.380 5.330 17.550 5.500 ;
        RECT 17.880 5.330 18.050 5.500 ;
        RECT 15.380 4.830 15.550 5.000 ;
        RECT 15.880 4.830 16.050 5.000 ;
        RECT 16.380 4.830 16.550 5.000 ;
        RECT 16.880 4.830 17.050 5.000 ;
        RECT 17.380 4.830 17.550 5.000 ;
        RECT 17.880 4.830 18.050 5.000 ;
        RECT 15.380 4.330 15.550 4.500 ;
        RECT 15.880 4.330 16.050 4.500 ;
        RECT 16.380 4.330 16.550 4.500 ;
        RECT 16.880 4.330 17.050 4.500 ;
        RECT 17.380 4.330 17.550 4.500 ;
        RECT 17.880 4.330 18.050 4.500 ;
        RECT 15.380 3.830 15.550 4.000 ;
        RECT 15.880 3.830 16.050 4.000 ;
        RECT 16.380 3.830 16.550 4.000 ;
        RECT 16.880 3.830 17.050 4.000 ;
        RECT 17.380 3.830 17.550 4.000 ;
        RECT 17.880 3.830 18.050 4.000 ;
        RECT 15.380 3.330 15.550 3.500 ;
        RECT 15.880 3.330 16.050 3.500 ;
        RECT 16.380 3.330 16.550 3.500 ;
        RECT 16.880 3.330 17.050 3.500 ;
        RECT 17.380 3.330 17.550 3.500 ;
        RECT 17.880 3.330 18.050 3.500 ;
        RECT 22.080 5.830 22.250 6.000 ;
        RECT 22.580 5.830 22.750 6.000 ;
        RECT 23.080 5.830 23.250 6.000 ;
        RECT 23.580 5.830 23.750 6.000 ;
        RECT 24.080 5.830 24.250 6.000 ;
        RECT 24.580 5.830 24.750 6.000 ;
        RECT 22.080 5.330 22.250 5.500 ;
        RECT 22.580 5.330 22.750 5.500 ;
        RECT 23.080 5.330 23.250 5.500 ;
        RECT 23.580 5.330 23.750 5.500 ;
        RECT 24.080 5.330 24.250 5.500 ;
        RECT 24.580 5.330 24.750 5.500 ;
        RECT 22.080 4.830 22.250 5.000 ;
        RECT 22.580 4.830 22.750 5.000 ;
        RECT 23.080 4.830 23.250 5.000 ;
        RECT 23.580 4.830 23.750 5.000 ;
        RECT 24.080 4.830 24.250 5.000 ;
        RECT 24.580 4.830 24.750 5.000 ;
        RECT 22.080 4.330 22.250 4.500 ;
        RECT 22.580 4.330 22.750 4.500 ;
        RECT 23.080 4.330 23.250 4.500 ;
        RECT 23.580 4.330 23.750 4.500 ;
        RECT 24.080 4.330 24.250 4.500 ;
        RECT 24.580 4.330 24.750 4.500 ;
        RECT 22.080 3.830 22.250 4.000 ;
        RECT 22.580 3.830 22.750 4.000 ;
        RECT 23.080 3.830 23.250 4.000 ;
        RECT 23.580 3.830 23.750 4.000 ;
        RECT 24.080 3.830 24.250 4.000 ;
        RECT 24.580 3.830 24.750 4.000 ;
        RECT 22.080 3.330 22.250 3.500 ;
        RECT 22.580 3.330 22.750 3.500 ;
        RECT 23.080 3.330 23.250 3.500 ;
        RECT 23.580 3.330 23.750 3.500 ;
        RECT 24.080 3.330 24.250 3.500 ;
        RECT 24.580 3.330 24.750 3.500 ;
        RECT 28.780 5.830 28.950 6.000 ;
        RECT 29.280 5.830 29.450 6.000 ;
        RECT 29.780 5.830 29.950 6.000 ;
        RECT 30.280 5.830 30.450 6.000 ;
        RECT 30.780 5.830 30.950 6.000 ;
        RECT 31.280 5.830 31.450 6.000 ;
        RECT 28.780 5.330 28.950 5.500 ;
        RECT 29.280 5.330 29.450 5.500 ;
        RECT 29.780 5.330 29.950 5.500 ;
        RECT 30.280 5.330 30.450 5.500 ;
        RECT 30.780 5.330 30.950 5.500 ;
        RECT 31.280 5.330 31.450 5.500 ;
        RECT 28.780 4.830 28.950 5.000 ;
        RECT 29.280 4.830 29.450 5.000 ;
        RECT 29.780 4.830 29.950 5.000 ;
        RECT 30.280 4.830 30.450 5.000 ;
        RECT 30.780 4.830 30.950 5.000 ;
        RECT 31.280 4.830 31.450 5.000 ;
        RECT 28.780 4.330 28.950 4.500 ;
        RECT 29.280 4.330 29.450 4.500 ;
        RECT 29.780 4.330 29.950 4.500 ;
        RECT 30.280 4.330 30.450 4.500 ;
        RECT 30.780 4.330 30.950 4.500 ;
        RECT 31.280 4.330 31.450 4.500 ;
        RECT 28.780 3.830 28.950 4.000 ;
        RECT 29.280 3.830 29.450 4.000 ;
        RECT 29.780 3.830 29.950 4.000 ;
        RECT 30.280 3.830 30.450 4.000 ;
        RECT 30.780 3.830 30.950 4.000 ;
        RECT 31.280 3.830 31.450 4.000 ;
        RECT 28.780 3.330 28.950 3.500 ;
        RECT 29.280 3.330 29.450 3.500 ;
        RECT 29.780 3.330 29.950 3.500 ;
        RECT 30.280 3.330 30.450 3.500 ;
        RECT 30.780 3.330 30.950 3.500 ;
        RECT 31.280 3.330 31.450 3.500 ;
        RECT 35.480 5.830 35.650 6.000 ;
        RECT 35.980 5.830 36.150 6.000 ;
        RECT 36.480 5.830 36.650 6.000 ;
        RECT 36.980 5.830 37.150 6.000 ;
        RECT 37.480 5.830 37.650 6.000 ;
        RECT 37.980 5.830 38.150 6.000 ;
        RECT 35.480 5.330 35.650 5.500 ;
        RECT 35.980 5.330 36.150 5.500 ;
        RECT 36.480 5.330 36.650 5.500 ;
        RECT 36.980 5.330 37.150 5.500 ;
        RECT 37.480 5.330 37.650 5.500 ;
        RECT 37.980 5.330 38.150 5.500 ;
        RECT 35.480 4.830 35.650 5.000 ;
        RECT 35.980 4.830 36.150 5.000 ;
        RECT 36.480 4.830 36.650 5.000 ;
        RECT 36.980 4.830 37.150 5.000 ;
        RECT 37.480 4.830 37.650 5.000 ;
        RECT 37.980 4.830 38.150 5.000 ;
        RECT 35.480 4.330 35.650 4.500 ;
        RECT 35.980 4.330 36.150 4.500 ;
        RECT 36.480 4.330 36.650 4.500 ;
        RECT 36.980 4.330 37.150 4.500 ;
        RECT 37.480 4.330 37.650 4.500 ;
        RECT 37.980 4.330 38.150 4.500 ;
        RECT 35.480 3.830 35.650 4.000 ;
        RECT 35.980 3.830 36.150 4.000 ;
        RECT 36.480 3.830 36.650 4.000 ;
        RECT 36.980 3.830 37.150 4.000 ;
        RECT 37.480 3.830 37.650 4.000 ;
        RECT 37.980 3.830 38.150 4.000 ;
        RECT 35.480 3.330 35.650 3.500 ;
        RECT 35.980 3.330 36.150 3.500 ;
        RECT 36.480 3.330 36.650 3.500 ;
        RECT 36.980 3.330 37.150 3.500 ;
        RECT 37.480 3.330 37.650 3.500 ;
        RECT 37.980 3.330 38.150 3.500 ;
        RECT 42.180 5.830 42.350 6.000 ;
        RECT 42.680 5.830 42.850 6.000 ;
        RECT 43.180 5.830 43.350 6.000 ;
        RECT 43.680 5.830 43.850 6.000 ;
        RECT 44.180 5.830 44.350 6.000 ;
        RECT 44.680 5.830 44.850 6.000 ;
        RECT 42.180 5.330 42.350 5.500 ;
        RECT 42.680 5.330 42.850 5.500 ;
        RECT 43.180 5.330 43.350 5.500 ;
        RECT 43.680 5.330 43.850 5.500 ;
        RECT 44.180 5.330 44.350 5.500 ;
        RECT 44.680 5.330 44.850 5.500 ;
        RECT 42.180 4.830 42.350 5.000 ;
        RECT 42.680 4.830 42.850 5.000 ;
        RECT 43.180 4.830 43.350 5.000 ;
        RECT 43.680 4.830 43.850 5.000 ;
        RECT 44.180 4.830 44.350 5.000 ;
        RECT 44.680 4.830 44.850 5.000 ;
        RECT 42.180 4.330 42.350 4.500 ;
        RECT 42.680 4.330 42.850 4.500 ;
        RECT 43.180 4.330 43.350 4.500 ;
        RECT 43.680 4.330 43.850 4.500 ;
        RECT 44.180 4.330 44.350 4.500 ;
        RECT 44.680 4.330 44.850 4.500 ;
        RECT 42.180 3.830 42.350 4.000 ;
        RECT 42.680 3.830 42.850 4.000 ;
        RECT 43.180 3.830 43.350 4.000 ;
        RECT 43.680 3.830 43.850 4.000 ;
        RECT 44.180 3.830 44.350 4.000 ;
        RECT 44.680 3.830 44.850 4.000 ;
        RECT 42.180 3.330 42.350 3.500 ;
        RECT 42.680 3.330 42.850 3.500 ;
        RECT 43.180 3.330 43.350 3.500 ;
        RECT 43.680 3.330 43.850 3.500 ;
        RECT 44.180 3.330 44.350 3.500 ;
        RECT 44.680 3.330 44.850 3.500 ;
        RECT 48.880 5.830 49.050 6.000 ;
        RECT 49.380 5.830 49.550 6.000 ;
        RECT 49.880 5.830 50.050 6.000 ;
        RECT 50.380 5.830 50.550 6.000 ;
        RECT 50.880 5.830 51.050 6.000 ;
        RECT 51.380 5.830 51.550 6.000 ;
        RECT 48.880 5.330 49.050 5.500 ;
        RECT 49.380 5.330 49.550 5.500 ;
        RECT 49.880 5.330 50.050 5.500 ;
        RECT 50.380 5.330 50.550 5.500 ;
        RECT 50.880 5.330 51.050 5.500 ;
        RECT 51.380 5.330 51.550 5.500 ;
        RECT 48.880 4.830 49.050 5.000 ;
        RECT 49.380 4.830 49.550 5.000 ;
        RECT 49.880 4.830 50.050 5.000 ;
        RECT 50.380 4.830 50.550 5.000 ;
        RECT 50.880 4.830 51.050 5.000 ;
        RECT 51.380 4.830 51.550 5.000 ;
        RECT 48.880 4.330 49.050 4.500 ;
        RECT 49.380 4.330 49.550 4.500 ;
        RECT 49.880 4.330 50.050 4.500 ;
        RECT 50.380 4.330 50.550 4.500 ;
        RECT 50.880 4.330 51.050 4.500 ;
        RECT 51.380 4.330 51.550 4.500 ;
        RECT 48.880 3.830 49.050 4.000 ;
        RECT 49.380 3.830 49.550 4.000 ;
        RECT 49.880 3.830 50.050 4.000 ;
        RECT 50.380 3.830 50.550 4.000 ;
        RECT 50.880 3.830 51.050 4.000 ;
        RECT 51.380 3.830 51.550 4.000 ;
        RECT 48.880 3.330 49.050 3.500 ;
        RECT 49.380 3.330 49.550 3.500 ;
        RECT 49.880 3.330 50.050 3.500 ;
        RECT 50.380 3.330 50.550 3.500 ;
        RECT 50.880 3.330 51.050 3.500 ;
        RECT 51.380 3.330 51.550 3.500 ;
      LAYER met1 ;
        RECT 1.820 3.170 51.780 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 51.264000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 6.745 5.755 7.105 ;
        RECT 0.945 2.655 1.305 6.745 ;
        RECT 5.395 2.655 5.755 6.745 ;
        RECT 0.945 2.295 5.755 2.655 ;
        RECT 7.645 6.745 12.455 7.105 ;
        RECT 7.645 2.655 8.005 6.745 ;
        RECT 12.095 2.655 12.455 6.745 ;
        RECT 7.645 2.295 12.455 2.655 ;
        RECT 14.345 6.745 19.155 7.105 ;
        RECT 14.345 2.655 14.705 6.745 ;
        RECT 18.795 2.655 19.155 6.745 ;
        RECT 14.345 2.295 19.155 2.655 ;
        RECT 21.045 6.745 25.855 7.105 ;
        RECT 21.045 2.655 21.405 6.745 ;
        RECT 25.495 2.655 25.855 6.745 ;
        RECT 21.045 2.295 25.855 2.655 ;
        RECT 27.745 6.745 32.555 7.105 ;
        RECT 27.745 2.655 28.105 6.745 ;
        RECT 32.195 2.655 32.555 6.745 ;
        RECT 27.745 2.295 32.555 2.655 ;
        RECT 34.445 6.745 39.255 7.105 ;
        RECT 34.445 2.655 34.805 6.745 ;
        RECT 38.895 2.655 39.255 6.745 ;
        RECT 34.445 2.295 39.255 2.655 ;
        RECT 41.145 6.745 45.955 7.105 ;
        RECT 41.145 2.655 41.505 6.745 ;
        RECT 45.595 2.655 45.955 6.745 ;
        RECT 41.145 2.295 45.955 2.655 ;
        RECT 47.845 6.745 52.655 7.105 ;
        RECT 47.845 2.655 48.205 6.745 ;
        RECT 52.295 2.655 52.655 6.745 ;
        RECT 47.845 2.295 52.655 2.655 ;
      LAYER mcon ;
        RECT 1.050 6.850 1.220 7.020 ;
        RECT 1.500 6.850 1.670 7.020 ;
        RECT 1.950 6.850 2.120 7.020 ;
        RECT 2.400 6.850 2.570 7.020 ;
        RECT 2.850 6.850 3.020 7.020 ;
        RECT 3.300 6.850 3.470 7.020 ;
        RECT 3.750 6.850 3.920 7.020 ;
        RECT 4.200 6.850 4.370 7.020 ;
        RECT 4.650 6.850 4.820 7.020 ;
        RECT 5.100 6.850 5.270 7.020 ;
        RECT 5.550 6.850 5.720 7.020 ;
        RECT 7.750 6.850 7.920 7.020 ;
        RECT 8.200 6.850 8.370 7.020 ;
        RECT 8.650 6.850 8.820 7.020 ;
        RECT 9.100 6.850 9.270 7.020 ;
        RECT 9.550 6.850 9.720 7.020 ;
        RECT 10.000 6.850 10.170 7.020 ;
        RECT 10.450 6.850 10.620 7.020 ;
        RECT 10.900 6.850 11.070 7.020 ;
        RECT 11.350 6.850 11.520 7.020 ;
        RECT 11.800 6.850 11.970 7.020 ;
        RECT 12.250 6.850 12.420 7.020 ;
        RECT 14.450 6.850 14.620 7.020 ;
        RECT 14.900 6.850 15.070 7.020 ;
        RECT 15.350 6.850 15.520 7.020 ;
        RECT 15.800 6.850 15.970 7.020 ;
        RECT 16.250 6.850 16.420 7.020 ;
        RECT 16.700 6.850 16.870 7.020 ;
        RECT 17.150 6.850 17.320 7.020 ;
        RECT 17.600 6.850 17.770 7.020 ;
        RECT 18.050 6.850 18.220 7.020 ;
        RECT 18.500 6.850 18.670 7.020 ;
        RECT 18.950 6.850 19.120 7.020 ;
        RECT 21.150 6.850 21.320 7.020 ;
        RECT 21.600 6.850 21.770 7.020 ;
        RECT 22.050 6.850 22.220 7.020 ;
        RECT 22.500 6.850 22.670 7.020 ;
        RECT 22.950 6.850 23.120 7.020 ;
        RECT 23.400 6.850 23.570 7.020 ;
        RECT 23.850 6.850 24.020 7.020 ;
        RECT 24.300 6.850 24.470 7.020 ;
        RECT 24.750 6.850 24.920 7.020 ;
        RECT 25.200 6.850 25.370 7.020 ;
        RECT 25.650 6.850 25.820 7.020 ;
        RECT 27.850 6.850 28.020 7.020 ;
        RECT 28.300 6.850 28.470 7.020 ;
        RECT 28.750 6.850 28.920 7.020 ;
        RECT 29.200 6.850 29.370 7.020 ;
        RECT 29.650 6.850 29.820 7.020 ;
        RECT 30.100 6.850 30.270 7.020 ;
        RECT 30.550 6.850 30.720 7.020 ;
        RECT 31.000 6.850 31.170 7.020 ;
        RECT 31.450 6.850 31.620 7.020 ;
        RECT 31.900 6.850 32.070 7.020 ;
        RECT 32.350 6.850 32.520 7.020 ;
        RECT 34.550 6.850 34.720 7.020 ;
        RECT 35.000 6.850 35.170 7.020 ;
        RECT 35.450 6.850 35.620 7.020 ;
        RECT 35.900 6.850 36.070 7.020 ;
        RECT 36.350 6.850 36.520 7.020 ;
        RECT 36.800 6.850 36.970 7.020 ;
        RECT 37.250 6.850 37.420 7.020 ;
        RECT 37.700 6.850 37.870 7.020 ;
        RECT 38.150 6.850 38.320 7.020 ;
        RECT 38.600 6.850 38.770 7.020 ;
        RECT 39.050 6.850 39.220 7.020 ;
        RECT 41.250 6.850 41.420 7.020 ;
        RECT 41.700 6.850 41.870 7.020 ;
        RECT 42.150 6.850 42.320 7.020 ;
        RECT 42.600 6.850 42.770 7.020 ;
        RECT 43.050 6.850 43.220 7.020 ;
        RECT 43.500 6.850 43.670 7.020 ;
        RECT 43.950 6.850 44.120 7.020 ;
        RECT 44.400 6.850 44.570 7.020 ;
        RECT 44.850 6.850 45.020 7.020 ;
        RECT 45.300 6.850 45.470 7.020 ;
        RECT 45.750 6.850 45.920 7.020 ;
        RECT 47.950 6.850 48.120 7.020 ;
        RECT 48.400 6.850 48.570 7.020 ;
        RECT 48.850 6.850 49.020 7.020 ;
        RECT 49.300 6.850 49.470 7.020 ;
        RECT 49.750 6.850 49.920 7.020 ;
        RECT 50.200 6.850 50.370 7.020 ;
        RECT 50.650 6.850 50.820 7.020 ;
        RECT 51.100 6.850 51.270 7.020 ;
        RECT 51.550 6.850 51.720 7.020 ;
        RECT 52.000 6.850 52.170 7.020 ;
        RECT 52.450 6.850 52.620 7.020 ;
      LAYER met1 ;
        RECT 0.950 6.750 52.650 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 107.630394 ;
    PORT
      LAYER pwell ;
        RECT 0.000 7.285 53.600 8.050 ;
        RECT 0.000 2.115 0.765 7.285 ;
        RECT 5.935 2.115 7.465 7.285 ;
        RECT 12.635 2.115 14.165 7.285 ;
        RECT 19.335 2.115 20.865 7.285 ;
        RECT 26.035 2.115 27.565 7.285 ;
        RECT 32.735 2.115 34.265 7.285 ;
        RECT 39.435 2.115 40.965 7.285 ;
        RECT 46.135 2.115 47.665 7.285 ;
        RECT 52.835 2.115 53.600 7.285 ;
        RECT 0.000 1.350 53.600 2.115 ;
      LAYER li1 ;
        RECT 0.130 7.425 53.470 7.920 ;
        RECT 0.130 1.975 0.625 7.425 ;
        RECT 6.075 1.975 7.325 7.425 ;
        RECT 12.775 1.975 14.025 7.425 ;
        RECT 19.475 1.975 20.725 7.425 ;
        RECT 26.175 1.975 27.425 7.425 ;
        RECT 32.875 1.975 34.125 7.425 ;
        RECT 39.575 1.975 40.825 7.425 ;
        RECT 46.275 1.975 47.525 7.425 ;
        RECT 52.975 1.975 53.470 7.425 ;
        RECT 0.130 1.480 53.470 1.975 ;
      LAYER mcon ;
        RECT 0.230 7.650 0.400 7.820 ;
        RECT 0.680 7.650 0.850 7.820 ;
        RECT 1.130 7.650 1.300 7.820 ;
        RECT 1.580 7.650 1.750 7.820 ;
        RECT 2.030 7.650 2.200 7.820 ;
        RECT 2.480 7.650 2.650 7.820 ;
        RECT 2.930 7.650 3.100 7.820 ;
        RECT 3.380 7.650 3.550 7.820 ;
        RECT 3.830 7.650 4.000 7.820 ;
        RECT 4.280 7.650 4.450 7.820 ;
        RECT 4.730 7.650 4.900 7.820 ;
        RECT 5.180 7.650 5.350 7.820 ;
        RECT 5.630 7.650 5.800 7.820 ;
        RECT 6.080 7.650 6.250 7.820 ;
        RECT 6.930 7.650 7.100 7.820 ;
        RECT 7.380 7.650 7.550 7.820 ;
        RECT 7.830 7.650 8.000 7.820 ;
        RECT 8.280 7.650 8.450 7.820 ;
        RECT 8.730 7.650 8.900 7.820 ;
        RECT 9.180 7.650 9.350 7.820 ;
        RECT 9.630 7.650 9.800 7.820 ;
        RECT 10.080 7.650 10.250 7.820 ;
        RECT 10.530 7.650 10.700 7.820 ;
        RECT 10.980 7.650 11.150 7.820 ;
        RECT 11.430 7.650 11.600 7.820 ;
        RECT 11.880 7.650 12.050 7.820 ;
        RECT 12.330 7.650 12.500 7.820 ;
        RECT 12.780 7.650 12.950 7.820 ;
        RECT 13.630 7.650 13.800 7.820 ;
        RECT 14.080 7.650 14.250 7.820 ;
        RECT 14.530 7.650 14.700 7.820 ;
        RECT 14.980 7.650 15.150 7.820 ;
        RECT 15.430 7.650 15.600 7.820 ;
        RECT 15.880 7.650 16.050 7.820 ;
        RECT 16.330 7.650 16.500 7.820 ;
        RECT 16.780 7.650 16.950 7.820 ;
        RECT 17.230 7.650 17.400 7.820 ;
        RECT 17.680 7.650 17.850 7.820 ;
        RECT 18.130 7.650 18.300 7.820 ;
        RECT 18.580 7.650 18.750 7.820 ;
        RECT 19.030 7.650 19.200 7.820 ;
        RECT 19.480 7.650 19.650 7.820 ;
        RECT 20.330 7.650 20.500 7.820 ;
        RECT 20.780 7.650 20.950 7.820 ;
        RECT 21.230 7.650 21.400 7.820 ;
        RECT 21.680 7.650 21.850 7.820 ;
        RECT 22.130 7.650 22.300 7.820 ;
        RECT 22.580 7.650 22.750 7.820 ;
        RECT 23.030 7.650 23.200 7.820 ;
        RECT 23.480 7.650 23.650 7.820 ;
        RECT 23.930 7.650 24.100 7.820 ;
        RECT 24.380 7.650 24.550 7.820 ;
        RECT 24.830 7.650 25.000 7.820 ;
        RECT 25.280 7.650 25.450 7.820 ;
        RECT 25.730 7.650 25.900 7.820 ;
        RECT 26.180 7.650 26.350 7.820 ;
        RECT 27.030 7.650 27.200 7.820 ;
        RECT 27.480 7.650 27.650 7.820 ;
        RECT 27.930 7.650 28.100 7.820 ;
        RECT 28.380 7.650 28.550 7.820 ;
        RECT 28.830 7.650 29.000 7.820 ;
        RECT 29.280 7.650 29.450 7.820 ;
        RECT 29.730 7.650 29.900 7.820 ;
        RECT 30.180 7.650 30.350 7.820 ;
        RECT 30.630 7.650 30.800 7.820 ;
        RECT 31.080 7.650 31.250 7.820 ;
        RECT 31.530 7.650 31.700 7.820 ;
        RECT 31.980 7.650 32.150 7.820 ;
        RECT 32.430 7.650 32.600 7.820 ;
        RECT 32.880 7.650 33.050 7.820 ;
        RECT 33.730 7.650 33.900 7.820 ;
        RECT 34.180 7.650 34.350 7.820 ;
        RECT 34.630 7.650 34.800 7.820 ;
        RECT 35.080 7.650 35.250 7.820 ;
        RECT 35.530 7.650 35.700 7.820 ;
        RECT 35.980 7.650 36.150 7.820 ;
        RECT 36.430 7.650 36.600 7.820 ;
        RECT 36.880 7.650 37.050 7.820 ;
        RECT 37.330 7.650 37.500 7.820 ;
        RECT 37.780 7.650 37.950 7.820 ;
        RECT 38.230 7.650 38.400 7.820 ;
        RECT 38.680 7.650 38.850 7.820 ;
        RECT 39.130 7.650 39.300 7.820 ;
        RECT 39.580 7.650 39.750 7.820 ;
        RECT 40.430 7.650 40.600 7.820 ;
        RECT 40.880 7.650 41.050 7.820 ;
        RECT 41.330 7.650 41.500 7.820 ;
        RECT 41.780 7.650 41.950 7.820 ;
        RECT 42.230 7.650 42.400 7.820 ;
        RECT 42.680 7.650 42.850 7.820 ;
        RECT 43.130 7.650 43.300 7.820 ;
        RECT 43.580 7.650 43.750 7.820 ;
        RECT 44.030 7.650 44.200 7.820 ;
        RECT 44.480 7.650 44.650 7.820 ;
        RECT 44.930 7.650 45.100 7.820 ;
        RECT 45.380 7.650 45.550 7.820 ;
        RECT 45.830 7.650 46.000 7.820 ;
        RECT 46.280 7.650 46.450 7.820 ;
        RECT 47.130 7.650 47.300 7.820 ;
        RECT 47.580 7.650 47.750 7.820 ;
        RECT 48.030 7.650 48.200 7.820 ;
        RECT 48.480 7.650 48.650 7.820 ;
        RECT 48.930 7.650 49.100 7.820 ;
        RECT 49.380 7.650 49.550 7.820 ;
        RECT 49.830 7.650 50.000 7.820 ;
        RECT 50.280 7.650 50.450 7.820 ;
        RECT 50.730 7.650 50.900 7.820 ;
        RECT 51.180 7.650 51.350 7.820 ;
        RECT 51.630 7.650 51.800 7.820 ;
        RECT 52.080 7.650 52.250 7.820 ;
        RECT 52.530 7.650 52.700 7.820 ;
        RECT 52.980 7.650 53.150 7.820 ;
      LAYER met1 ;
        RECT 0.130 7.500 53.470 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 53.600 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 1.850 9.250 2.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 3.850 9.250 4.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 5.850 9.250 6.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 7.850 9.250 8.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 9.850 9.250 10.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 11.850 9.250 12.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 13.850 9.250 14.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 15.850 9.250 16.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 17.850 9.250 18.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
        RECT 19.850 9.250 20.150 9.550 ;
        RECT 20.850 9.250 21.150 9.550 ;
        RECT 21.850 9.250 22.150 9.550 ;
        RECT 22.850 9.250 23.150 9.550 ;
        RECT 23.850 9.250 24.150 9.550 ;
        RECT 24.850 9.250 25.150 9.550 ;
        RECT 25.850 9.250 26.150 9.550 ;
        RECT 26.850 9.250 27.150 9.550 ;
        RECT 27.850 9.250 28.150 9.550 ;
        RECT 28.850 9.250 29.150 9.550 ;
        RECT 29.850 9.250 30.150 9.550 ;
        RECT 30.850 9.250 31.150 9.550 ;
        RECT 31.850 9.250 32.150 9.550 ;
        RECT 32.850 9.250 33.150 9.550 ;
        RECT 33.850 9.250 34.150 9.550 ;
        RECT 34.850 9.250 35.150 9.550 ;
        RECT 35.850 9.250 36.150 9.550 ;
        RECT 36.850 9.250 37.150 9.550 ;
        RECT 37.850 9.250 38.150 9.550 ;
        RECT 38.850 9.250 39.150 9.550 ;
        RECT 39.850 9.250 40.150 9.550 ;
        RECT 40.850 9.250 41.150 9.550 ;
        RECT 41.850 9.250 42.150 9.550 ;
        RECT 42.850 9.250 43.150 9.550 ;
        RECT 43.850 9.250 44.150 9.550 ;
        RECT 44.850 9.250 45.150 9.550 ;
        RECT 45.850 9.250 46.150 9.550 ;
        RECT 46.850 9.250 47.150 9.550 ;
        RECT 47.850 9.250 48.150 9.550 ;
        RECT 48.850 9.250 49.150 9.550 ;
        RECT 49.850 9.250 50.150 9.550 ;
        RECT 50.850 9.250 51.150 9.550 ;
        RECT 51.850 9.250 52.150 9.550 ;
        RECT 52.850 9.250 53.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 53.600 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 53.600 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.850 -0.150 21.150 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.850 -0.150 23.150 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.850 -0.150 25.150 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.850 -0.150 27.150 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.850 -0.150 29.150 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.850 -0.150 31.150 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.850 -0.150 33.150 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.850 -0.150 35.150 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.850 -0.150 37.150 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.850 -0.150 39.150 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.850 -0.150 41.150 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.850 -0.150 43.150 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.850 -0.150 45.150 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
        RECT 46.850 -0.150 47.150 0.150 ;
        RECT 47.850 -0.150 48.150 0.150 ;
        RECT 48.850 -0.150 49.150 0.150 ;
        RECT 49.850 -0.150 50.150 0.150 ;
        RECT 50.850 -0.150 51.150 0.150 ;
        RECT 51.850 -0.150 52.150 0.150 ;
        RECT 52.850 -0.150 53.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 53.600 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_8

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.070 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.890 0.720 3.070 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.490 8.450 3.070 8.750 ;
        RECT 2.835 7.020 3.005 8.450 ;
        RECT 2.835 6.930 3.010 7.020 ;
        RECT 2.840 2.980 3.010 6.930 ;
      LAYER mcon ;
        RECT 2.840 3.060 3.010 6.940 ;
      LAYER met1 ;
        RECT 2.810 3.000 3.040 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.550 3.270 0.720 7.020 ;
        RECT 0.545 2.980 0.720 3.270 ;
        RECT 0.545 2.150 0.715 2.980 ;
        RECT 0.490 1.850 3.070 2.150 ;
      LAYER mcon ;
        RECT 0.550 3.060 0.720 6.940 ;
      LAYER met1 ;
        RECT 0.520 3.000 0.750 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 3.070 9.550 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 3.070 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.100 0.150 3.170 7.130 ;
      LAYER li1 ;
        RECT 0.140 0.150 0.440 1.200 ;
        RECT 0.000 -0.150 3.070 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 3.070 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.430 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 3.430 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 3.430 8.950 ;
        RECT 3.015 8.245 3.185 8.650 ;
        RECT 3.015 8.130 3.190 8.245 ;
        RECT 3.020 1.755 3.190 8.130 ;
      LAYER mcon ;
        RECT 3.020 1.835 3.190 8.165 ;
      LAYER met1 ;
        RECT 2.990 1.775 3.220 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.730 1.870 0.900 8.245 ;
        RECT 0.725 1.755 0.900 1.870 ;
        RECT 0.725 1.350 0.895 1.755 ;
        RECT 0.490 1.050 3.430 1.350 ;
      LAYER mcon ;
        RECT 0.730 1.835 0.900 8.165 ;
      LAYER met1 ;
        RECT 0.700 1.775 0.930 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.100 1.470 3.530 9.700 ;
        RECT 0.490 1.465 3.430 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 3.430 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 3.430 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 3.430 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 3.430 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_res_xhigh_po_2p85_1
  CLASS CORE ;
  FOREIGN sky130_asc_res_xhigh_po_2p85_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.200 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.000 5.375 2.160 8.225 ;
      LAYER mcon ;
        RECT 0.090 5.455 2.075 8.145 ;
      LAYER met1 ;
        RECT 0.055 5.395 2.105 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.575 2.160 3.425 ;
      LAYER mcon ;
        RECT 0.090 0.655 2.075 3.345 ;
      LAYER met1 ;
        RECT 0.055 0.595 2.105 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 12.200 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 1.850 9.250 2.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 3.850 9.250 4.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 5.850 9.250 6.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 7.850 9.250 8.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 9.850 9.250 10.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 12.200 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.300 12.200 8.250 ;
      LAYER li1 ;
        RECT 4.560 0.150 7.640 4.850 ;
        RECT 0.000 -0.150 12.200 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 12.200 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 10.040 0.575 12.200 8.225 ;
      LAYER mcon ;
        RECT 10.125 5.455 12.110 8.145 ;
        RECT 10.125 0.655 12.110 3.345 ;
      LAYER met1 ;
        RECT 10.095 5.395 12.145 8.205 ;
        RECT 10.040 0.575 12.200 5.395 ;
  END
END sky130_asc_res_xhigh_po_2p85_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.535 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 138.530 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 138.530 8.950 ;
        RECT 3.015 1.755 3.185 8.650 ;
        RECT 7.595 1.755 7.765 8.650 ;
        RECT 12.175 1.755 12.345 8.650 ;
        RECT 16.755 1.755 16.925 8.650 ;
        RECT 21.335 1.755 21.505 8.650 ;
        RECT 25.915 1.755 26.085 8.650 ;
        RECT 30.495 1.755 30.665 8.650 ;
        RECT 35.075 1.755 35.245 8.650 ;
        RECT 39.655 1.755 39.825 8.650 ;
        RECT 44.235 1.755 44.405 8.650 ;
        RECT 48.815 1.755 48.985 8.650 ;
        RECT 53.395 1.755 53.565 8.650 ;
        RECT 57.975 1.755 58.145 8.650 ;
        RECT 62.555 1.755 62.725 8.650 ;
        RECT 67.135 1.755 67.305 8.650 ;
        RECT 71.715 1.755 71.885 8.650 ;
        RECT 76.295 1.755 76.465 8.650 ;
        RECT 80.875 1.755 81.045 8.650 ;
        RECT 85.455 1.755 85.625 8.650 ;
        RECT 90.035 1.755 90.205 8.650 ;
        RECT 94.615 1.755 94.785 8.650 ;
        RECT 99.195 1.755 99.365 8.650 ;
        RECT 103.775 1.755 103.945 8.650 ;
        RECT 108.355 1.755 108.525 8.650 ;
        RECT 112.935 1.755 113.105 8.650 ;
        RECT 117.515 1.755 117.685 8.650 ;
        RECT 122.095 1.755 122.265 8.650 ;
        RECT 126.675 1.755 126.845 8.650 ;
        RECT 131.255 1.755 131.425 8.650 ;
        RECT 135.835 1.755 136.005 8.650 ;
      LAYER mcon ;
        RECT 3.015 1.835 3.185 8.165 ;
        RECT 7.595 1.835 7.765 8.165 ;
        RECT 12.175 1.835 12.345 8.165 ;
        RECT 16.755 1.835 16.925 8.165 ;
        RECT 21.335 1.835 21.505 8.165 ;
        RECT 25.915 1.835 26.085 8.165 ;
        RECT 30.495 1.835 30.665 8.165 ;
        RECT 35.075 1.835 35.245 8.165 ;
        RECT 39.655 1.835 39.825 8.165 ;
        RECT 44.235 1.835 44.405 8.165 ;
        RECT 48.815 1.835 48.985 8.165 ;
        RECT 53.395 1.835 53.565 8.165 ;
        RECT 57.975 1.835 58.145 8.165 ;
        RECT 62.555 1.835 62.725 8.165 ;
        RECT 67.135 1.835 67.305 8.165 ;
        RECT 71.715 1.835 71.885 8.165 ;
        RECT 76.295 1.835 76.465 8.165 ;
        RECT 80.875 1.835 81.045 8.165 ;
        RECT 85.455 1.835 85.625 8.165 ;
        RECT 90.035 1.835 90.205 8.165 ;
        RECT 94.615 1.835 94.785 8.165 ;
        RECT 99.195 1.835 99.365 8.165 ;
        RECT 103.775 1.835 103.945 8.165 ;
        RECT 108.355 1.835 108.525 8.165 ;
        RECT 112.935 1.835 113.105 8.165 ;
        RECT 117.515 1.835 117.685 8.165 ;
        RECT 122.095 1.835 122.265 8.165 ;
        RECT 126.675 1.835 126.845 8.165 ;
        RECT 131.255 1.835 131.425 8.165 ;
        RECT 135.835 1.835 136.005 8.165 ;
      LAYER met1 ;
        RECT 2.985 1.775 3.215 8.225 ;
        RECT 7.565 1.775 7.795 8.225 ;
        RECT 12.145 1.775 12.375 8.225 ;
        RECT 16.725 1.775 16.955 8.225 ;
        RECT 21.305 1.775 21.535 8.225 ;
        RECT 25.885 1.775 26.115 8.225 ;
        RECT 30.465 1.775 30.695 8.225 ;
        RECT 35.045 1.775 35.275 8.225 ;
        RECT 39.625 1.775 39.855 8.225 ;
        RECT 44.205 1.775 44.435 8.225 ;
        RECT 48.785 1.775 49.015 8.225 ;
        RECT 53.365 1.775 53.595 8.225 ;
        RECT 57.945 1.775 58.175 8.225 ;
        RECT 62.525 1.775 62.755 8.225 ;
        RECT 67.105 1.775 67.335 8.225 ;
        RECT 71.685 1.775 71.915 8.225 ;
        RECT 76.265 1.775 76.495 8.225 ;
        RECT 80.845 1.775 81.075 8.225 ;
        RECT 85.425 1.775 85.655 8.225 ;
        RECT 90.005 1.775 90.235 8.225 ;
        RECT 94.585 1.775 94.815 8.225 ;
        RECT 99.165 1.775 99.395 8.225 ;
        RECT 103.745 1.775 103.975 8.225 ;
        RECT 108.325 1.775 108.555 8.225 ;
        RECT 112.905 1.775 113.135 8.225 ;
        RECT 117.485 1.775 117.715 8.225 ;
        RECT 122.065 1.775 122.295 8.225 ;
        RECT 126.645 1.775 126.875 8.225 ;
        RECT 131.225 1.775 131.455 8.225 ;
        RECT 135.805 1.775 136.035 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.350 0.895 8.245 ;
        RECT 5.305 1.350 5.475 8.245 ;
        RECT 9.885 1.350 10.055 8.245 ;
        RECT 14.465 1.350 14.635 8.245 ;
        RECT 19.045 1.350 19.215 8.245 ;
        RECT 23.625 1.350 23.795 8.245 ;
        RECT 28.205 1.350 28.375 8.245 ;
        RECT 32.785 1.350 32.955 8.245 ;
        RECT 37.365 1.350 37.535 8.245 ;
        RECT 41.945 1.350 42.115 8.245 ;
        RECT 46.525 1.350 46.695 8.245 ;
        RECT 51.105 1.350 51.275 8.245 ;
        RECT 55.685 1.350 55.855 8.245 ;
        RECT 60.265 1.350 60.435 8.245 ;
        RECT 64.845 1.350 65.015 8.245 ;
        RECT 69.425 1.350 69.595 8.245 ;
        RECT 74.005 1.350 74.175 8.245 ;
        RECT 78.585 1.350 78.755 8.245 ;
        RECT 83.165 1.350 83.335 8.245 ;
        RECT 87.745 1.350 87.915 8.245 ;
        RECT 92.325 1.350 92.495 8.245 ;
        RECT 96.905 1.350 97.075 8.245 ;
        RECT 101.485 1.350 101.655 8.245 ;
        RECT 106.065 1.350 106.235 8.245 ;
        RECT 110.645 1.350 110.815 8.245 ;
        RECT 115.225 1.350 115.395 8.245 ;
        RECT 119.805 1.350 119.975 8.245 ;
        RECT 124.385 1.350 124.555 8.245 ;
        RECT 128.965 1.350 129.135 8.245 ;
        RECT 133.545 1.350 133.715 8.245 ;
        RECT 138.125 1.350 138.295 8.245 ;
        RECT 0.490 1.050 138.530 1.350 ;
      LAYER mcon ;
        RECT 0.725 1.835 0.895 8.165 ;
        RECT 5.305 1.835 5.475 8.165 ;
        RECT 9.885 1.835 10.055 8.165 ;
        RECT 14.465 1.835 14.635 8.165 ;
        RECT 19.045 1.835 19.215 8.165 ;
        RECT 23.625 1.835 23.795 8.165 ;
        RECT 28.205 1.835 28.375 8.165 ;
        RECT 32.785 1.835 32.955 8.165 ;
        RECT 37.365 1.835 37.535 8.165 ;
        RECT 41.945 1.835 42.115 8.165 ;
        RECT 46.525 1.835 46.695 8.165 ;
        RECT 51.105 1.835 51.275 8.165 ;
        RECT 55.685 1.835 55.855 8.165 ;
        RECT 60.265 1.835 60.435 8.165 ;
        RECT 64.845 1.835 65.015 8.165 ;
        RECT 69.425 1.835 69.595 8.165 ;
        RECT 74.005 1.835 74.175 8.165 ;
        RECT 78.585 1.835 78.755 8.165 ;
        RECT 83.165 1.835 83.335 8.165 ;
        RECT 87.745 1.835 87.915 8.165 ;
        RECT 92.325 1.835 92.495 8.165 ;
        RECT 96.905 1.835 97.075 8.165 ;
        RECT 101.485 1.835 101.655 8.165 ;
        RECT 106.065 1.835 106.235 8.165 ;
        RECT 110.645 1.835 110.815 8.165 ;
        RECT 115.225 1.835 115.395 8.165 ;
        RECT 119.805 1.835 119.975 8.165 ;
        RECT 124.385 1.835 124.555 8.165 ;
        RECT 128.965 1.835 129.135 8.165 ;
        RECT 133.545 1.835 133.715 8.165 ;
        RECT 138.125 1.835 138.295 8.165 ;
      LAYER met1 ;
        RECT 0.695 1.775 0.925 8.225 ;
        RECT 5.275 1.775 5.505 8.225 ;
        RECT 9.855 1.775 10.085 8.225 ;
        RECT 14.435 1.775 14.665 8.225 ;
        RECT 19.015 1.775 19.245 8.225 ;
        RECT 23.595 1.775 23.825 8.225 ;
        RECT 28.175 1.775 28.405 8.225 ;
        RECT 32.755 1.775 32.985 8.225 ;
        RECT 37.335 1.775 37.565 8.225 ;
        RECT 41.915 1.775 42.145 8.225 ;
        RECT 46.495 1.775 46.725 8.225 ;
        RECT 51.075 1.775 51.305 8.225 ;
        RECT 55.655 1.775 55.885 8.225 ;
        RECT 60.235 1.775 60.465 8.225 ;
        RECT 64.815 1.775 65.045 8.225 ;
        RECT 69.395 1.775 69.625 8.225 ;
        RECT 73.975 1.775 74.205 8.225 ;
        RECT 78.555 1.775 78.785 8.225 ;
        RECT 83.135 1.775 83.365 8.225 ;
        RECT 87.715 1.775 87.945 8.225 ;
        RECT 92.295 1.775 92.525 8.225 ;
        RECT 96.875 1.775 97.105 8.225 ;
        RECT 101.455 1.775 101.685 8.225 ;
        RECT 106.035 1.775 106.265 8.225 ;
        RECT 110.615 1.775 110.845 8.225 ;
        RECT 115.195 1.775 115.425 8.225 ;
        RECT 119.775 1.775 120.005 8.225 ;
        RECT 124.355 1.775 124.585 8.225 ;
        RECT 128.935 1.775 129.165 8.225 ;
        RECT 133.515 1.775 133.745 8.225 ;
        RECT 138.095 1.775 138.325 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 8.535 138.530 9.700 ;
        RECT 0.000 1.470 138.535 8.535 ;
        RECT 0.485 1.465 138.535 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 138.530 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
        RECT 15.340 9.250 15.640 9.550 ;
        RECT 17.340 9.250 17.640 9.550 ;
        RECT 19.340 9.250 19.640 9.550 ;
        RECT 21.340 9.250 21.640 9.550 ;
        RECT 23.340 9.250 23.640 9.550 ;
        RECT 25.340 9.250 25.640 9.550 ;
        RECT 27.340 9.250 27.640 9.550 ;
        RECT 29.340 9.250 29.640 9.550 ;
        RECT 31.340 9.250 31.640 9.550 ;
        RECT 33.340 9.250 33.640 9.550 ;
        RECT 35.340 9.250 35.640 9.550 ;
        RECT 37.340 9.250 37.640 9.550 ;
        RECT 39.340 9.250 39.640 9.550 ;
        RECT 41.340 9.250 41.640 9.550 ;
        RECT 43.340 9.250 43.640 9.550 ;
        RECT 45.340 9.250 45.640 9.550 ;
        RECT 47.340 9.250 47.640 9.550 ;
        RECT 49.340 9.250 49.640 9.550 ;
        RECT 51.340 9.250 51.640 9.550 ;
        RECT 53.340 9.250 53.640 9.550 ;
        RECT 55.340 9.250 55.640 9.550 ;
        RECT 57.340 9.250 57.640 9.550 ;
        RECT 59.340 9.250 59.640 9.550 ;
        RECT 61.340 9.250 61.640 9.550 ;
        RECT 63.340 9.250 63.640 9.550 ;
        RECT 65.340 9.250 65.640 9.550 ;
        RECT 67.340 9.250 67.640 9.550 ;
        RECT 69.340 9.250 69.640 9.550 ;
        RECT 71.340 9.250 71.640 9.550 ;
        RECT 73.340 9.250 73.640 9.550 ;
        RECT 75.340 9.250 75.640 9.550 ;
        RECT 77.340 9.250 77.640 9.550 ;
        RECT 79.340 9.250 79.640 9.550 ;
        RECT 81.340 9.250 81.640 9.550 ;
        RECT 83.340 9.250 83.640 9.550 ;
        RECT 85.340 9.250 85.640 9.550 ;
        RECT 87.340 9.250 87.640 9.550 ;
        RECT 89.340 9.250 89.640 9.550 ;
        RECT 91.340 9.250 91.640 9.550 ;
        RECT 93.340 9.250 93.640 9.550 ;
        RECT 95.340 9.250 95.640 9.550 ;
        RECT 97.340 9.250 97.640 9.550 ;
        RECT 99.340 9.250 99.640 9.550 ;
        RECT 101.340 9.250 101.640 9.550 ;
        RECT 103.340 9.250 103.640 9.550 ;
        RECT 105.340 9.250 105.640 9.550 ;
        RECT 107.340 9.250 107.640 9.550 ;
        RECT 109.340 9.250 109.640 9.550 ;
        RECT 111.340 9.250 111.640 9.550 ;
        RECT 113.340 9.250 113.640 9.550 ;
        RECT 115.340 9.250 115.640 9.550 ;
        RECT 117.340 9.250 117.640 9.550 ;
        RECT 119.340 9.250 119.640 9.550 ;
        RECT 121.340 9.250 121.640 9.550 ;
        RECT 123.340 9.250 123.640 9.550 ;
        RECT 125.340 9.250 125.640 9.550 ;
        RECT 127.340 9.250 127.640 9.550 ;
        RECT 129.340 9.250 129.640 9.550 ;
        RECT 131.340 9.250 131.640 9.550 ;
        RECT 133.340 9.250 133.640 9.550 ;
        RECT 135.340 9.250 135.640 9.550 ;
        RECT 137.340 9.250 137.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 138.530 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 138.530 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
        RECT 15.340 -0.150 15.640 0.150 ;
        RECT 17.340 -0.150 17.640 0.150 ;
        RECT 19.340 -0.150 19.640 0.150 ;
        RECT 21.340 -0.150 21.640 0.150 ;
        RECT 23.340 -0.150 23.640 0.150 ;
        RECT 25.340 -0.150 25.640 0.150 ;
        RECT 27.340 -0.150 27.640 0.150 ;
        RECT 29.340 -0.150 29.640 0.150 ;
        RECT 31.340 -0.150 31.640 0.150 ;
        RECT 33.340 -0.150 33.640 0.150 ;
        RECT 35.340 -0.150 35.640 0.150 ;
        RECT 37.340 -0.150 37.640 0.150 ;
        RECT 39.340 -0.150 39.640 0.150 ;
        RECT 41.340 -0.150 41.640 0.150 ;
        RECT 43.340 -0.150 43.640 0.150 ;
        RECT 45.340 -0.150 45.640 0.150 ;
        RECT 47.340 -0.150 47.640 0.150 ;
        RECT 49.340 -0.150 49.640 0.150 ;
        RECT 51.340 -0.150 51.640 0.150 ;
        RECT 53.340 -0.150 53.640 0.150 ;
        RECT 55.340 -0.150 55.640 0.150 ;
        RECT 57.340 -0.150 57.640 0.150 ;
        RECT 59.340 -0.150 59.640 0.150 ;
        RECT 61.340 -0.150 61.640 0.150 ;
        RECT 63.340 -0.150 63.640 0.150 ;
        RECT 65.340 -0.150 65.640 0.150 ;
        RECT 67.340 -0.150 67.640 0.150 ;
        RECT 69.340 -0.150 69.640 0.150 ;
        RECT 71.340 -0.150 71.640 0.150 ;
        RECT 73.340 -0.150 73.640 0.150 ;
        RECT 75.340 -0.150 75.640 0.150 ;
        RECT 77.340 -0.150 77.640 0.150 ;
        RECT 79.340 -0.150 79.640 0.150 ;
        RECT 81.340 -0.150 81.640 0.150 ;
        RECT 83.340 -0.150 83.640 0.150 ;
        RECT 85.340 -0.150 85.640 0.150 ;
        RECT 87.340 -0.150 87.640 0.150 ;
        RECT 89.340 -0.150 89.640 0.150 ;
        RECT 91.340 -0.150 91.640 0.150 ;
        RECT 93.340 -0.150 93.640 0.150 ;
        RECT 95.340 -0.150 95.640 0.150 ;
        RECT 97.340 -0.150 97.640 0.150 ;
        RECT 99.340 -0.150 99.640 0.150 ;
        RECT 101.340 -0.150 101.640 0.150 ;
        RECT 103.340 -0.150 103.640 0.150 ;
        RECT 105.340 -0.150 105.640 0.150 ;
        RECT 107.340 -0.150 107.640 0.150 ;
        RECT 109.340 -0.150 109.640 0.150 ;
        RECT 111.340 -0.150 111.640 0.150 ;
        RECT 113.340 -0.150 113.640 0.150 ;
        RECT 115.340 -0.150 115.640 0.150 ;
        RECT 117.340 -0.150 117.640 0.150 ;
        RECT 119.340 -0.150 119.640 0.150 ;
        RECT 121.340 -0.150 121.640 0.150 ;
        RECT 123.340 -0.150 123.640 0.150 ;
        RECT 125.340 -0.150 125.640 0.150 ;
        RECT 127.340 -0.150 127.640 0.150 ;
        RECT 129.340 -0.150 129.640 0.150 ;
        RECT 131.340 -0.150 131.640 0.150 ;
        RECT 133.340 -0.150 133.640 0.150 ;
        RECT 135.340 -0.150 135.640 0.150 ;
        RECT 137.340 -0.150 137.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 138.530 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60

#--------EOF---------

MACRO sky130_asc_res_xhigh_po_2p85_2
  CLASS CORE ;
  FOREIGN sky130_asc_res_xhigh_po_2p85_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.070 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.005 5.375 2.165 8.225 ;
      LAYER mcon ;
        RECT 0.095 5.455 2.080 8.145 ;
      LAYER met1 ;
        RECT 0.060 5.395 2.110 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.005 0.575 2.165 3.425 ;
      LAYER mcon ;
        RECT 0.095 0.655 2.080 3.345 ;
      LAYER met1 ;
        RECT 0.060 0.595 2.110 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 9.250 15.070 9.550 ;
      LAYER mcon ;
        RECT 0.860 9.250 1.160 9.550 ;
        RECT 1.860 9.250 2.160 9.550 ;
        RECT 2.860 9.250 3.160 9.550 ;
        RECT 3.860 9.250 4.160 9.550 ;
        RECT 4.860 9.250 5.160 9.550 ;
        RECT 5.860 9.250 6.160 9.550 ;
        RECT 6.860 9.250 7.160 9.550 ;
        RECT 7.860 9.250 8.160 9.550 ;
        RECT 8.860 9.250 9.160 9.550 ;
        RECT 9.860 9.250 10.160 9.550 ;
        RECT 10.860 9.250 11.160 9.550 ;
        RECT 11.860 9.250 12.160 9.550 ;
        RECT 12.860 9.250 13.160 9.550 ;
        RECT 13.860 9.250 14.160 9.550 ;
      LAYER met1 ;
        RECT 0.010 9.100 15.070 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.440 -0.300 13.640 8.250 ;
      LAYER li1 ;
        RECT 6.000 0.150 9.080 4.850 ;
        RECT 0.010 -0.150 15.070 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 1.860 -0.150 2.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 3.860 -0.150 4.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 5.860 -0.150 6.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 7.860 -0.150 8.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 9.860 -0.150 10.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 11.860 -0.150 12.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
        RECT 13.860 -0.150 14.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 15.070 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 12.915 0.575 15.075 8.225 ;
      LAYER mcon ;
        RECT 13.000 5.455 14.985 8.145 ;
        RECT 13.000 0.655 14.985 3.345 ;
      LAYER met1 ;
        RECT 12.970 5.395 15.020 8.205 ;
        RECT 12.915 0.575 15.075 5.395 ;
  END
END sky130_asc_res_xhigh_po_2p85_2

#--------EOF---------

MACRO sky130_asc_pnp_05v5_W3p40L3p40_1
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.700 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.559999 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.965 5.085 6.435 ;
      LAYER mcon ;
        RECT 1.980 5.830 2.150 6.000 ;
        RECT 2.480 5.830 2.650 6.000 ;
        RECT 2.980 5.830 3.150 6.000 ;
        RECT 3.480 5.830 3.650 6.000 ;
        RECT 3.980 5.830 4.150 6.000 ;
        RECT 4.480 5.830 4.650 6.000 ;
        RECT 1.980 5.330 2.150 5.500 ;
        RECT 2.480 5.330 2.650 5.500 ;
        RECT 2.980 5.330 3.150 5.500 ;
        RECT 3.480 5.330 3.650 5.500 ;
        RECT 3.980 5.330 4.150 5.500 ;
        RECT 4.480 5.330 4.650 5.500 ;
        RECT 1.980 4.830 2.150 5.000 ;
        RECT 2.480 4.830 2.650 5.000 ;
        RECT 2.980 4.830 3.150 5.000 ;
        RECT 3.480 4.830 3.650 5.000 ;
        RECT 3.980 4.830 4.150 5.000 ;
        RECT 4.480 4.830 4.650 5.000 ;
        RECT 1.980 4.330 2.150 4.500 ;
        RECT 2.480 4.330 2.650 4.500 ;
        RECT 2.980 4.330 3.150 4.500 ;
        RECT 3.480 4.330 3.650 4.500 ;
        RECT 3.980 4.330 4.150 4.500 ;
        RECT 4.480 4.330 4.650 4.500 ;
        RECT 1.980 3.830 2.150 4.000 ;
        RECT 2.480 3.830 2.650 4.000 ;
        RECT 2.980 3.830 3.150 4.000 ;
        RECT 3.480 3.830 3.650 4.000 ;
        RECT 3.980 3.830 4.150 4.000 ;
        RECT 4.480 3.830 4.650 4.000 ;
        RECT 1.980 3.330 2.150 3.500 ;
        RECT 2.480 3.330 2.650 3.500 ;
        RECT 2.980 3.330 3.150 3.500 ;
        RECT 3.480 3.330 3.650 3.500 ;
        RECT 3.980 3.330 4.150 3.500 ;
        RECT 4.480 3.330 4.650 3.500 ;
      LAYER met1 ;
        RECT 1.825 3.175 4.875 6.225 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 6.408000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 6.745 5.755 7.105 ;
        RECT 0.945 2.655 1.305 6.745 ;
        RECT 5.395 2.655 5.755 6.745 ;
        RECT 0.945 2.295 5.755 2.655 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.988700 ;
    PORT
      LAYER pwell ;
        RECT 0.000 7.285 6.700 8.050 ;
        RECT 0.000 2.115 0.765 7.285 ;
        RECT 5.935 2.115 6.700 7.285 ;
        RECT 0.000 1.350 6.700 2.115 ;
      LAYER li1 ;
        RECT 0.130 7.425 6.570 7.920 ;
        RECT 0.130 1.975 0.625 7.425 ;
        RECT 6.075 1.975 6.570 7.425 ;
        RECT 0.130 1.480 6.570 1.975 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 6.700 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 1.850 9.250 2.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 3.850 9.250 4.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 5.850 9.250 6.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 6.700 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 6.700 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 6.700 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_12
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.615 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 154.800003 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 28.610 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.223000 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 28.610 8.950 ;
        RECT 3.015 1.755 3.185 8.650 ;
        RECT 7.595 1.755 7.765 8.650 ;
        RECT 12.175 1.755 12.345 8.650 ;
        RECT 16.755 1.755 16.925 8.650 ;
        RECT 21.335 1.755 21.505 8.650 ;
        RECT 25.915 1.755 26.085 8.650 ;
      LAYER mcon ;
        RECT 3.015 1.835 3.185 8.165 ;
        RECT 7.595 1.835 7.765 8.165 ;
        RECT 12.175 1.835 12.345 8.165 ;
        RECT 16.755 1.835 16.925 8.165 ;
        RECT 21.335 1.835 21.505 8.165 ;
        RECT 25.915 1.835 26.085 8.165 ;
      LAYER met1 ;
        RECT 2.985 1.775 3.215 8.225 ;
        RECT 7.565 1.775 7.795 8.225 ;
        RECT 12.145 1.775 12.375 8.225 ;
        RECT 16.725 1.775 16.955 8.225 ;
        RECT 21.305 1.775 21.535 8.225 ;
        RECT 25.885 1.775 26.115 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.093500 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.350 0.895 8.245 ;
        RECT 5.305 1.350 5.475 8.245 ;
        RECT 9.885 1.350 10.055 8.245 ;
        RECT 14.465 1.350 14.635 8.245 ;
        RECT 19.045 1.350 19.215 8.245 ;
        RECT 23.625 1.350 23.795 8.245 ;
        RECT 28.205 1.350 28.375 8.245 ;
        RECT 0.490 1.050 28.610 1.350 ;
      LAYER mcon ;
        RECT 0.725 1.835 0.895 8.165 ;
        RECT 5.305 1.835 5.475 8.165 ;
        RECT 9.885 1.835 10.055 8.165 ;
        RECT 14.465 1.835 14.635 8.165 ;
        RECT 19.045 1.835 19.215 8.165 ;
        RECT 23.625 1.835 23.795 8.165 ;
        RECT 28.205 1.835 28.375 8.165 ;
      LAYER met1 ;
        RECT 0.695 1.775 0.925 8.225 ;
        RECT 5.275 1.775 5.505 8.225 ;
        RECT 9.855 1.775 10.085 8.225 ;
        RECT 14.435 1.775 14.665 8.225 ;
        RECT 19.015 1.775 19.245 8.225 ;
        RECT 23.595 1.775 23.825 8.225 ;
        RECT 28.175 1.775 28.405 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 8.535 28.610 9.700 ;
        RECT 0.000 1.470 28.615 8.535 ;
        RECT 0.485 1.465 28.615 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 28.610 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
        RECT 15.340 9.250 15.640 9.550 ;
        RECT 17.340 9.250 17.640 9.550 ;
        RECT 19.340 9.250 19.640 9.550 ;
        RECT 21.340 9.250 21.640 9.550 ;
        RECT 23.340 9.250 23.640 9.550 ;
        RECT 25.340 9.250 25.640 9.550 ;
        RECT 27.340 9.250 27.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 28.610 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 28.610 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
        RECT 15.340 -0.150 15.640 0.150 ;
        RECT 17.340 -0.150 17.640 0.150 ;
        RECT 19.340 -0.150 19.640 0.150 ;
        RECT 21.340 -0.150 21.640 0.150 ;
        RECT 23.340 -0.150 23.640 0.150 ;
        RECT 25.340 -0.150 25.640 0.150 ;
        RECT 27.340 -0.150 27.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 28.610 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_12

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.875 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 14.870 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 14.870 8.950 ;
        RECT 3.015 1.755 3.185 8.650 ;
        RECT 7.595 1.755 7.765 8.650 ;
        RECT 12.175 1.755 12.345 8.650 ;
      LAYER mcon ;
        RECT 3.015 1.835 3.185 8.165 ;
        RECT 7.595 1.835 7.765 8.165 ;
        RECT 12.175 1.835 12.345 8.165 ;
      LAYER met1 ;
        RECT 2.985 1.775 3.215 8.225 ;
        RECT 7.565 1.775 7.795 8.225 ;
        RECT 12.145 1.775 12.375 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.350 0.895 8.245 ;
        RECT 5.305 1.350 5.475 8.245 ;
        RECT 9.885 1.350 10.055 8.245 ;
        RECT 14.465 1.350 14.635 8.245 ;
        RECT 0.490 1.050 14.870 1.350 ;
      LAYER mcon ;
        RECT 0.725 1.835 0.895 8.165 ;
        RECT 5.305 1.835 5.475 8.165 ;
        RECT 9.885 1.835 10.055 8.165 ;
        RECT 14.465 1.835 14.635 8.165 ;
      LAYER met1 ;
        RECT 0.695 1.775 0.925 8.225 ;
        RECT 5.275 1.775 5.505 8.225 ;
        RECT 9.855 1.775 10.085 8.225 ;
        RECT 14.435 1.775 14.665 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 8.535 14.870 9.700 ;
        RECT 0.000 1.470 14.875 8.535 ;
        RECT 0.485 1.465 14.875 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 14.870 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 14.870 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 14.870 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 14.870 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_6

#--------EOF---------

MACRO sky130_asc_pnp_05v5_W3p40L3p40_7
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_7 ;
  ORIGIN 0.000 0.000 ;
  SIZE 46.900 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 80.919998 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.965 5.085 6.435 ;
        RECT 8.315 2.965 11.785 6.435 ;
        RECT 15.015 2.965 18.485 6.435 ;
        RECT 21.715 2.965 25.185 6.435 ;
        RECT 28.415 2.965 31.885 6.435 ;
        RECT 35.115 2.965 38.585 6.435 ;
        RECT 41.815 2.965 45.285 6.435 ;
      LAYER mcon ;
        RECT 1.980 5.830 2.150 6.000 ;
        RECT 2.480 5.830 2.650 6.000 ;
        RECT 2.980 5.830 3.150 6.000 ;
        RECT 3.480 5.830 3.650 6.000 ;
        RECT 3.980 5.830 4.150 6.000 ;
        RECT 4.480 5.830 4.650 6.000 ;
        RECT 1.980 5.330 2.150 5.500 ;
        RECT 2.480 5.330 2.650 5.500 ;
        RECT 2.980 5.330 3.150 5.500 ;
        RECT 3.480 5.330 3.650 5.500 ;
        RECT 3.980 5.330 4.150 5.500 ;
        RECT 4.480 5.330 4.650 5.500 ;
        RECT 1.980 4.830 2.150 5.000 ;
        RECT 2.480 4.830 2.650 5.000 ;
        RECT 2.980 4.830 3.150 5.000 ;
        RECT 3.480 4.830 3.650 5.000 ;
        RECT 3.980 4.830 4.150 5.000 ;
        RECT 4.480 4.830 4.650 5.000 ;
        RECT 1.980 4.330 2.150 4.500 ;
        RECT 2.480 4.330 2.650 4.500 ;
        RECT 2.980 4.330 3.150 4.500 ;
        RECT 3.480 4.330 3.650 4.500 ;
        RECT 3.980 4.330 4.150 4.500 ;
        RECT 4.480 4.330 4.650 4.500 ;
        RECT 1.980 3.830 2.150 4.000 ;
        RECT 2.480 3.830 2.650 4.000 ;
        RECT 2.980 3.830 3.150 4.000 ;
        RECT 3.480 3.830 3.650 4.000 ;
        RECT 3.980 3.830 4.150 4.000 ;
        RECT 4.480 3.830 4.650 4.000 ;
        RECT 1.980 3.330 2.150 3.500 ;
        RECT 2.480 3.330 2.650 3.500 ;
        RECT 2.980 3.330 3.150 3.500 ;
        RECT 3.480 3.330 3.650 3.500 ;
        RECT 3.980 3.330 4.150 3.500 ;
        RECT 4.480 3.330 4.650 3.500 ;
        RECT 8.680 5.830 8.850 6.000 ;
        RECT 9.180 5.830 9.350 6.000 ;
        RECT 9.680 5.830 9.850 6.000 ;
        RECT 10.180 5.830 10.350 6.000 ;
        RECT 10.680 5.830 10.850 6.000 ;
        RECT 11.180 5.830 11.350 6.000 ;
        RECT 8.680 5.330 8.850 5.500 ;
        RECT 9.180 5.330 9.350 5.500 ;
        RECT 9.680 5.330 9.850 5.500 ;
        RECT 10.180 5.330 10.350 5.500 ;
        RECT 10.680 5.330 10.850 5.500 ;
        RECT 11.180 5.330 11.350 5.500 ;
        RECT 8.680 4.830 8.850 5.000 ;
        RECT 9.180 4.830 9.350 5.000 ;
        RECT 9.680 4.830 9.850 5.000 ;
        RECT 10.180 4.830 10.350 5.000 ;
        RECT 10.680 4.830 10.850 5.000 ;
        RECT 11.180 4.830 11.350 5.000 ;
        RECT 8.680 4.330 8.850 4.500 ;
        RECT 9.180 4.330 9.350 4.500 ;
        RECT 9.680 4.330 9.850 4.500 ;
        RECT 10.180 4.330 10.350 4.500 ;
        RECT 10.680 4.330 10.850 4.500 ;
        RECT 11.180 4.330 11.350 4.500 ;
        RECT 8.680 3.830 8.850 4.000 ;
        RECT 9.180 3.830 9.350 4.000 ;
        RECT 9.680 3.830 9.850 4.000 ;
        RECT 10.180 3.830 10.350 4.000 ;
        RECT 10.680 3.830 10.850 4.000 ;
        RECT 11.180 3.830 11.350 4.000 ;
        RECT 8.680 3.330 8.850 3.500 ;
        RECT 9.180 3.330 9.350 3.500 ;
        RECT 9.680 3.330 9.850 3.500 ;
        RECT 10.180 3.330 10.350 3.500 ;
        RECT 10.680 3.330 10.850 3.500 ;
        RECT 11.180 3.330 11.350 3.500 ;
        RECT 15.380 5.830 15.550 6.000 ;
        RECT 15.880 5.830 16.050 6.000 ;
        RECT 16.380 5.830 16.550 6.000 ;
        RECT 16.880 5.830 17.050 6.000 ;
        RECT 17.380 5.830 17.550 6.000 ;
        RECT 17.880 5.830 18.050 6.000 ;
        RECT 15.380 5.330 15.550 5.500 ;
        RECT 15.880 5.330 16.050 5.500 ;
        RECT 16.380 5.330 16.550 5.500 ;
        RECT 16.880 5.330 17.050 5.500 ;
        RECT 17.380 5.330 17.550 5.500 ;
        RECT 17.880 5.330 18.050 5.500 ;
        RECT 15.380 4.830 15.550 5.000 ;
        RECT 15.880 4.830 16.050 5.000 ;
        RECT 16.380 4.830 16.550 5.000 ;
        RECT 16.880 4.830 17.050 5.000 ;
        RECT 17.380 4.830 17.550 5.000 ;
        RECT 17.880 4.830 18.050 5.000 ;
        RECT 15.380 4.330 15.550 4.500 ;
        RECT 15.880 4.330 16.050 4.500 ;
        RECT 16.380 4.330 16.550 4.500 ;
        RECT 16.880 4.330 17.050 4.500 ;
        RECT 17.380 4.330 17.550 4.500 ;
        RECT 17.880 4.330 18.050 4.500 ;
        RECT 15.380 3.830 15.550 4.000 ;
        RECT 15.880 3.830 16.050 4.000 ;
        RECT 16.380 3.830 16.550 4.000 ;
        RECT 16.880 3.830 17.050 4.000 ;
        RECT 17.380 3.830 17.550 4.000 ;
        RECT 17.880 3.830 18.050 4.000 ;
        RECT 15.380 3.330 15.550 3.500 ;
        RECT 15.880 3.330 16.050 3.500 ;
        RECT 16.380 3.330 16.550 3.500 ;
        RECT 16.880 3.330 17.050 3.500 ;
        RECT 17.380 3.330 17.550 3.500 ;
        RECT 17.880 3.330 18.050 3.500 ;
        RECT 22.080 5.830 22.250 6.000 ;
        RECT 22.580 5.830 22.750 6.000 ;
        RECT 23.080 5.830 23.250 6.000 ;
        RECT 23.580 5.830 23.750 6.000 ;
        RECT 24.080 5.830 24.250 6.000 ;
        RECT 24.580 5.830 24.750 6.000 ;
        RECT 22.080 5.330 22.250 5.500 ;
        RECT 22.580 5.330 22.750 5.500 ;
        RECT 23.080 5.330 23.250 5.500 ;
        RECT 23.580 5.330 23.750 5.500 ;
        RECT 24.080 5.330 24.250 5.500 ;
        RECT 24.580 5.330 24.750 5.500 ;
        RECT 22.080 4.830 22.250 5.000 ;
        RECT 22.580 4.830 22.750 5.000 ;
        RECT 23.080 4.830 23.250 5.000 ;
        RECT 23.580 4.830 23.750 5.000 ;
        RECT 24.080 4.830 24.250 5.000 ;
        RECT 24.580 4.830 24.750 5.000 ;
        RECT 22.080 4.330 22.250 4.500 ;
        RECT 22.580 4.330 22.750 4.500 ;
        RECT 23.080 4.330 23.250 4.500 ;
        RECT 23.580 4.330 23.750 4.500 ;
        RECT 24.080 4.330 24.250 4.500 ;
        RECT 24.580 4.330 24.750 4.500 ;
        RECT 22.080 3.830 22.250 4.000 ;
        RECT 22.580 3.830 22.750 4.000 ;
        RECT 23.080 3.830 23.250 4.000 ;
        RECT 23.580 3.830 23.750 4.000 ;
        RECT 24.080 3.830 24.250 4.000 ;
        RECT 24.580 3.830 24.750 4.000 ;
        RECT 22.080 3.330 22.250 3.500 ;
        RECT 22.580 3.330 22.750 3.500 ;
        RECT 23.080 3.330 23.250 3.500 ;
        RECT 23.580 3.330 23.750 3.500 ;
        RECT 24.080 3.330 24.250 3.500 ;
        RECT 24.580 3.330 24.750 3.500 ;
        RECT 28.780 5.830 28.950 6.000 ;
        RECT 29.280 5.830 29.450 6.000 ;
        RECT 29.780 5.830 29.950 6.000 ;
        RECT 30.280 5.830 30.450 6.000 ;
        RECT 30.780 5.830 30.950 6.000 ;
        RECT 31.280 5.830 31.450 6.000 ;
        RECT 28.780 5.330 28.950 5.500 ;
        RECT 29.280 5.330 29.450 5.500 ;
        RECT 29.780 5.330 29.950 5.500 ;
        RECT 30.280 5.330 30.450 5.500 ;
        RECT 30.780 5.330 30.950 5.500 ;
        RECT 31.280 5.330 31.450 5.500 ;
        RECT 28.780 4.830 28.950 5.000 ;
        RECT 29.280 4.830 29.450 5.000 ;
        RECT 29.780 4.830 29.950 5.000 ;
        RECT 30.280 4.830 30.450 5.000 ;
        RECT 30.780 4.830 30.950 5.000 ;
        RECT 31.280 4.830 31.450 5.000 ;
        RECT 28.780 4.330 28.950 4.500 ;
        RECT 29.280 4.330 29.450 4.500 ;
        RECT 29.780 4.330 29.950 4.500 ;
        RECT 30.280 4.330 30.450 4.500 ;
        RECT 30.780 4.330 30.950 4.500 ;
        RECT 31.280 4.330 31.450 4.500 ;
        RECT 28.780 3.830 28.950 4.000 ;
        RECT 29.280 3.830 29.450 4.000 ;
        RECT 29.780 3.830 29.950 4.000 ;
        RECT 30.280 3.830 30.450 4.000 ;
        RECT 30.780 3.830 30.950 4.000 ;
        RECT 31.280 3.830 31.450 4.000 ;
        RECT 28.780 3.330 28.950 3.500 ;
        RECT 29.280 3.330 29.450 3.500 ;
        RECT 29.780 3.330 29.950 3.500 ;
        RECT 30.280 3.330 30.450 3.500 ;
        RECT 30.780 3.330 30.950 3.500 ;
        RECT 31.280 3.330 31.450 3.500 ;
        RECT 35.480 5.830 35.650 6.000 ;
        RECT 35.980 5.830 36.150 6.000 ;
        RECT 36.480 5.830 36.650 6.000 ;
        RECT 36.980 5.830 37.150 6.000 ;
        RECT 37.480 5.830 37.650 6.000 ;
        RECT 37.980 5.830 38.150 6.000 ;
        RECT 35.480 5.330 35.650 5.500 ;
        RECT 35.980 5.330 36.150 5.500 ;
        RECT 36.480 5.330 36.650 5.500 ;
        RECT 36.980 5.330 37.150 5.500 ;
        RECT 37.480 5.330 37.650 5.500 ;
        RECT 37.980 5.330 38.150 5.500 ;
        RECT 35.480 4.830 35.650 5.000 ;
        RECT 35.980 4.830 36.150 5.000 ;
        RECT 36.480 4.830 36.650 5.000 ;
        RECT 36.980 4.830 37.150 5.000 ;
        RECT 37.480 4.830 37.650 5.000 ;
        RECT 37.980 4.830 38.150 5.000 ;
        RECT 35.480 4.330 35.650 4.500 ;
        RECT 35.980 4.330 36.150 4.500 ;
        RECT 36.480 4.330 36.650 4.500 ;
        RECT 36.980 4.330 37.150 4.500 ;
        RECT 37.480 4.330 37.650 4.500 ;
        RECT 37.980 4.330 38.150 4.500 ;
        RECT 35.480 3.830 35.650 4.000 ;
        RECT 35.980 3.830 36.150 4.000 ;
        RECT 36.480 3.830 36.650 4.000 ;
        RECT 36.980 3.830 37.150 4.000 ;
        RECT 37.480 3.830 37.650 4.000 ;
        RECT 37.980 3.830 38.150 4.000 ;
        RECT 35.480 3.330 35.650 3.500 ;
        RECT 35.980 3.330 36.150 3.500 ;
        RECT 36.480 3.330 36.650 3.500 ;
        RECT 36.980 3.330 37.150 3.500 ;
        RECT 37.480 3.330 37.650 3.500 ;
        RECT 37.980 3.330 38.150 3.500 ;
        RECT 42.180 5.830 42.350 6.000 ;
        RECT 42.680 5.830 42.850 6.000 ;
        RECT 43.180 5.830 43.350 6.000 ;
        RECT 43.680 5.830 43.850 6.000 ;
        RECT 44.180 5.830 44.350 6.000 ;
        RECT 44.680 5.830 44.850 6.000 ;
        RECT 42.180 5.330 42.350 5.500 ;
        RECT 42.680 5.330 42.850 5.500 ;
        RECT 43.180 5.330 43.350 5.500 ;
        RECT 43.680 5.330 43.850 5.500 ;
        RECT 44.180 5.330 44.350 5.500 ;
        RECT 44.680 5.330 44.850 5.500 ;
        RECT 42.180 4.830 42.350 5.000 ;
        RECT 42.680 4.830 42.850 5.000 ;
        RECT 43.180 4.830 43.350 5.000 ;
        RECT 43.680 4.830 43.850 5.000 ;
        RECT 44.180 4.830 44.350 5.000 ;
        RECT 44.680 4.830 44.850 5.000 ;
        RECT 42.180 4.330 42.350 4.500 ;
        RECT 42.680 4.330 42.850 4.500 ;
        RECT 43.180 4.330 43.350 4.500 ;
        RECT 43.680 4.330 43.850 4.500 ;
        RECT 44.180 4.330 44.350 4.500 ;
        RECT 44.680 4.330 44.850 4.500 ;
        RECT 42.180 3.830 42.350 4.000 ;
        RECT 42.680 3.830 42.850 4.000 ;
        RECT 43.180 3.830 43.350 4.000 ;
        RECT 43.680 3.830 43.850 4.000 ;
        RECT 44.180 3.830 44.350 4.000 ;
        RECT 44.680 3.830 44.850 4.000 ;
        RECT 42.180 3.330 42.350 3.500 ;
        RECT 42.680 3.330 42.850 3.500 ;
        RECT 43.180 3.330 43.350 3.500 ;
        RECT 43.680 3.330 43.850 3.500 ;
        RECT 44.180 3.330 44.350 3.500 ;
        RECT 44.680 3.330 44.850 3.500 ;
      LAYER met1 ;
        RECT 1.820 3.170 45.310 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 187.102295 ;
    ANTENNADIFFAREA 138.823303 ;
    PORT
      LAYER pwell ;
        RECT 0.000 7.285 46.900 8.050 ;
        RECT 0.000 2.115 0.765 7.285 ;
        RECT 5.935 2.115 7.465 7.285 ;
        RECT 12.635 2.115 14.165 7.285 ;
        RECT 19.335 2.115 20.865 7.285 ;
        RECT 26.035 2.115 27.565 7.285 ;
        RECT 32.735 2.115 34.265 7.285 ;
        RECT 39.435 2.115 40.965 7.285 ;
        RECT 46.135 2.115 46.900 7.285 ;
        RECT 0.000 1.350 46.900 2.115 ;
      LAYER li1 ;
        RECT 0.130 7.050 46.785 7.920 ;
        RECT 0.130 2.350 0.625 7.050 ;
        RECT 0.945 6.745 5.755 7.050 ;
        RECT 0.945 2.655 1.305 6.745 ;
        RECT 5.395 2.655 5.755 6.745 ;
        RECT 0.945 2.350 5.755 2.655 ;
        RECT 6.075 2.350 7.325 7.050 ;
        RECT 7.645 6.745 12.455 7.050 ;
        RECT 7.645 2.655 8.005 6.745 ;
        RECT 12.095 2.655 12.455 6.745 ;
        RECT 7.645 2.350 12.455 2.655 ;
        RECT 12.775 2.350 14.025 7.050 ;
        RECT 14.345 6.745 19.155 7.050 ;
        RECT 14.345 2.655 14.705 6.745 ;
        RECT 18.795 2.655 19.155 6.745 ;
        RECT 14.345 2.350 19.155 2.655 ;
        RECT 19.475 2.350 20.725 7.050 ;
        RECT 21.045 6.745 25.855 7.050 ;
        RECT 21.045 2.655 21.405 6.745 ;
        RECT 25.495 2.655 25.855 6.745 ;
        RECT 21.045 2.350 25.855 2.655 ;
        RECT 26.175 2.350 27.425 7.050 ;
        RECT 27.745 6.745 32.555 7.050 ;
        RECT 27.745 2.655 28.105 6.745 ;
        RECT 32.195 2.655 32.555 6.745 ;
        RECT 27.745 2.350 32.555 2.655 ;
        RECT 32.875 2.350 34.125 7.050 ;
        RECT 34.445 6.745 39.255 7.050 ;
        RECT 34.445 2.655 34.805 6.745 ;
        RECT 38.895 2.655 39.255 6.745 ;
        RECT 34.445 2.350 39.255 2.655 ;
        RECT 39.575 2.350 40.825 7.050 ;
        RECT 41.145 6.745 45.955 7.050 ;
        RECT 41.145 2.655 41.505 6.745 ;
        RECT 45.595 2.655 45.955 6.745 ;
        RECT 41.145 2.350 45.955 2.655 ;
        RECT 46.275 2.350 46.770 7.050 ;
        RECT 0.130 1.480 46.785 2.350 ;
    END
  END Base
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 46.900 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 1.850 9.250 2.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 3.850 9.250 4.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 5.850 9.250 6.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 7.850 9.250 8.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 9.850 9.250 10.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 11.850 9.250 12.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 13.850 9.250 14.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 15.850 9.250 16.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 17.850 9.250 18.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
        RECT 19.850 9.250 20.150 9.550 ;
        RECT 20.850 9.250 21.150 9.550 ;
        RECT 21.850 9.250 22.150 9.550 ;
        RECT 22.850 9.250 23.150 9.550 ;
        RECT 23.850 9.250 24.150 9.550 ;
        RECT 24.850 9.250 25.150 9.550 ;
        RECT 25.850 9.250 26.150 9.550 ;
        RECT 26.850 9.250 27.150 9.550 ;
        RECT 27.850 9.250 28.150 9.550 ;
        RECT 28.850 9.250 29.150 9.550 ;
        RECT 29.850 9.250 30.150 9.550 ;
        RECT 30.850 9.250 31.150 9.550 ;
        RECT 31.850 9.250 32.150 9.550 ;
        RECT 32.850 9.250 33.150 9.550 ;
        RECT 33.850 9.250 34.150 9.550 ;
        RECT 34.850 9.250 35.150 9.550 ;
        RECT 35.850 9.250 36.150 9.550 ;
        RECT 36.850 9.250 37.150 9.550 ;
        RECT 37.850 9.250 38.150 9.550 ;
        RECT 38.850 9.250 39.150 9.550 ;
        RECT 39.850 9.250 40.150 9.550 ;
        RECT 40.850 9.250 41.150 9.550 ;
        RECT 41.850 9.250 42.150 9.550 ;
        RECT 42.850 9.250 43.150 9.550 ;
        RECT 43.850 9.250 44.150 9.550 ;
        RECT 44.850 9.250 45.150 9.550 ;
        RECT 45.850 9.250 46.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 46.900 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 46.900 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.850 -0.150 21.150 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.850 -0.150 23.150 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.850 -0.150 25.150 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.850 -0.150 27.150 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.850 -0.150 29.150 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.850 -0.150 31.150 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.850 -0.150 33.150 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.850 -0.150 35.150 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.850 -0.150 37.150 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.850 -0.150 39.150 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.850 -0.150 41.150 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.850 -0.150 43.150 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.850 -0.150 45.150 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 46.900 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_7

#--------EOF---------

MACRO sky130_asc_cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_asc_cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.855 BY 9.400 ;
  SITE unitasc ;
  PIN Cin
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.250 35.850 8.450 ;
        RECT 0.000 5.250 35.855 8.250 ;
        RECT 0.000 4.750 35.850 5.250 ;
        RECT 0.000 1.750 35.855 4.750 ;
      LAYER via3 ;
        RECT 3.080 5.390 3.400 8.110 ;
        RECT 6.675 5.390 6.995 8.110 ;
        RECT 10.270 5.390 10.590 8.110 ;
        RECT 13.865 5.390 14.185 8.110 ;
        RECT 17.460 5.390 17.780 8.110 ;
        RECT 21.055 5.390 21.375 8.110 ;
        RECT 24.650 5.390 24.970 8.110 ;
        RECT 28.245 5.390 28.565 8.110 ;
        RECT 31.840 5.390 32.160 8.110 ;
        RECT 35.435 5.390 35.755 8.110 ;
        RECT 3.080 1.890 3.400 4.610 ;
        RECT 6.675 1.890 6.995 4.610 ;
        RECT 10.270 1.890 10.590 4.610 ;
        RECT 13.865 1.890 14.185 4.610 ;
        RECT 17.460 1.890 17.780 4.610 ;
        RECT 21.055 1.890 21.375 4.610 ;
        RECT 24.650 1.890 24.970 4.610 ;
        RECT 28.245 1.890 28.565 4.610 ;
        RECT 31.840 1.890 32.160 4.610 ;
        RECT 35.435 1.890 35.755 4.610 ;
      LAYER met4 ;
        RECT 3.000 5.310 3.480 8.190 ;
        RECT 6.595 5.310 7.075 8.190 ;
        RECT 10.190 5.310 10.670 8.190 ;
        RECT 13.785 5.310 14.265 8.190 ;
        RECT 17.380 5.310 17.860 8.190 ;
        RECT 20.975 5.310 21.455 8.190 ;
        RECT 24.570 5.310 25.050 8.190 ;
        RECT 28.165 5.310 28.645 8.190 ;
        RECT 31.760 5.310 32.240 8.190 ;
        RECT 35.355 5.310 35.835 8.190 ;
        RECT 3.000 1.810 3.480 4.690 ;
        RECT 6.595 1.810 7.075 4.690 ;
        RECT 10.190 1.810 10.670 4.690 ;
        RECT 13.785 1.810 14.265 4.690 ;
        RECT 17.380 1.810 17.860 4.690 ;
        RECT 20.975 1.810 21.455 4.690 ;
        RECT 24.570 1.810 25.050 4.690 ;
        RECT 28.165 1.810 28.645 4.690 ;
        RECT 31.760 1.810 32.240 4.690 ;
        RECT 35.355 1.810 35.835 4.690 ;
    END
  END Cin
  PIN Cout
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 0.700 7.555 2.300 7.650 ;
        RECT 4.300 7.555 5.900 7.650 ;
        RECT 7.900 7.555 9.500 7.650 ;
        RECT 11.500 7.555 13.100 7.650 ;
        RECT 15.100 7.555 16.700 7.650 ;
        RECT 18.700 7.555 20.300 7.650 ;
        RECT 22.300 7.555 23.900 7.650 ;
        RECT 25.900 7.555 27.500 7.650 ;
        RECT 29.500 7.555 31.100 7.650 ;
        RECT 33.100 7.555 34.700 7.650 ;
        RECT 0.700 5.945 2.310 7.555 ;
        RECT 4.295 5.945 5.905 7.555 ;
        RECT 7.890 5.945 9.500 7.555 ;
        RECT 11.485 5.945 13.100 7.555 ;
        RECT 15.080 5.945 16.700 7.555 ;
        RECT 18.675 5.945 20.300 7.555 ;
        RECT 22.270 5.945 23.900 7.555 ;
        RECT 25.865 5.945 27.500 7.555 ;
        RECT 29.460 5.945 31.100 7.555 ;
        RECT 33.055 5.945 34.700 7.555 ;
        RECT 0.700 4.055 2.300 5.945 ;
        RECT 4.300 4.055 5.900 5.945 ;
        RECT 7.900 4.055 9.500 5.945 ;
        RECT 11.500 4.055 13.100 5.945 ;
        RECT 15.100 4.055 16.700 5.945 ;
        RECT 18.700 4.055 20.300 5.945 ;
        RECT 22.300 4.055 23.900 5.945 ;
        RECT 25.900 4.055 27.500 5.945 ;
        RECT 29.500 4.055 31.100 5.945 ;
        RECT 33.100 4.055 34.700 5.945 ;
        RECT 0.700 2.445 2.310 4.055 ;
        RECT 4.295 2.445 5.905 4.055 ;
        RECT 7.890 2.445 9.500 4.055 ;
        RECT 11.485 2.445 13.100 4.055 ;
        RECT 15.080 2.445 16.700 4.055 ;
        RECT 18.675 2.445 20.300 4.055 ;
        RECT 22.270 2.445 23.900 4.055 ;
        RECT 25.865 2.445 27.500 4.055 ;
        RECT 29.460 2.445 31.100 4.055 ;
        RECT 33.055 2.445 34.700 4.055 ;
        RECT 0.700 1.450 2.300 2.445 ;
        RECT 4.300 1.450 5.900 2.445 ;
        RECT 7.900 1.450 9.500 2.445 ;
        RECT 11.500 1.450 13.100 2.445 ;
        RECT 15.100 1.450 16.700 2.445 ;
        RECT 18.700 1.450 20.300 2.445 ;
        RECT 22.300 1.450 23.900 2.445 ;
        RECT 25.900 1.450 27.500 2.445 ;
        RECT 29.500 1.450 31.100 2.445 ;
        RECT 33.100 1.450 34.700 2.445 ;
        RECT 0.010 0.950 35.850 1.450 ;
    END
  END Cout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 9.250 35.850 9.550 ;
      LAYER mcon ;
        RECT 0.860 9.250 1.160 9.550 ;
        RECT 2.860 9.250 3.160 9.550 ;
        RECT 4.860 9.250 5.160 9.550 ;
        RECT 6.860 9.250 7.160 9.550 ;
        RECT 8.860 9.250 9.160 9.550 ;
        RECT 10.860 9.250 11.160 9.550 ;
        RECT 12.860 9.250 13.160 9.550 ;
        RECT 14.860 9.250 15.160 9.550 ;
        RECT 16.860 9.250 17.160 9.550 ;
        RECT 18.860 9.250 19.160 9.550 ;
        RECT 20.860 9.250 21.160 9.550 ;
        RECT 22.860 9.250 23.160 9.550 ;
        RECT 24.860 9.250 25.160 9.550 ;
        RECT 26.860 9.250 27.160 9.550 ;
        RECT 28.860 9.250 29.160 9.550 ;
        RECT 30.860 9.250 31.160 9.550 ;
        RECT 32.860 9.250 33.160 9.550 ;
        RECT 34.860 9.250 35.160 9.550 ;
      LAYER met1 ;
        RECT 0.010 9.100 35.850 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.010 -0.150 35.850 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
        RECT 14.860 -0.150 15.160 0.150 ;
        RECT 16.860 -0.150 17.160 0.150 ;
        RECT 18.860 -0.150 19.160 0.150 ;
        RECT 20.860 -0.150 21.160 0.150 ;
        RECT 22.860 -0.150 23.160 0.150 ;
        RECT 24.860 -0.150 25.160 0.150 ;
        RECT 26.860 -0.150 27.160 0.150 ;
        RECT 28.860 -0.150 29.160 0.150 ;
        RECT 30.860 -0.150 31.160 0.150 ;
        RECT 32.860 -0.150 33.160 0.150 ;
        RECT 34.860 -0.150 35.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 35.850 0.300 ;
    END
  END VGND
END sky130_asc_cap_mim_m3_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.750 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 21.750 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 21.750 8.950 ;
        RECT 3.015 8.245 3.185 8.650 ;
        RECT 7.595 8.245 7.765 8.650 ;
        RECT 12.175 8.245 12.345 8.650 ;
        RECT 16.755 8.245 16.925 8.650 ;
        RECT 21.335 8.245 21.505 8.650 ;
        RECT 3.015 8.130 3.190 8.245 ;
        RECT 7.595 8.130 7.770 8.245 ;
        RECT 12.175 8.130 12.350 8.245 ;
        RECT 16.755 8.130 16.930 8.245 ;
        RECT 21.335 8.130 21.510 8.245 ;
        RECT 3.020 1.755 3.190 8.130 ;
        RECT 7.600 1.755 7.770 8.130 ;
        RECT 12.180 1.755 12.350 8.130 ;
        RECT 16.760 1.755 16.930 8.130 ;
        RECT 21.340 1.755 21.510 8.130 ;
      LAYER mcon ;
        RECT 3.020 1.835 3.190 8.165 ;
        RECT 7.600 1.835 7.770 8.165 ;
        RECT 12.180 1.835 12.350 8.165 ;
        RECT 16.760 1.835 16.930 8.165 ;
        RECT 21.340 1.835 21.510 8.165 ;
      LAYER met1 ;
        RECT 2.990 1.775 3.220 8.225 ;
        RECT 7.570 1.775 7.800 8.225 ;
        RECT 12.150 1.775 12.380 8.225 ;
        RECT 16.730 1.775 16.960 8.225 ;
        RECT 21.310 1.775 21.540 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.730 1.870 0.900 8.245 ;
        RECT 5.310 1.870 5.480 8.245 ;
        RECT 9.890 1.870 10.060 8.245 ;
        RECT 14.470 1.870 14.640 8.245 ;
        RECT 19.050 1.870 19.220 8.245 ;
        RECT 0.725 1.755 0.900 1.870 ;
        RECT 5.305 1.755 5.480 1.870 ;
        RECT 9.885 1.755 10.060 1.870 ;
        RECT 14.465 1.755 14.640 1.870 ;
        RECT 19.045 1.755 19.220 1.870 ;
        RECT 0.725 1.350 0.895 1.755 ;
        RECT 5.305 1.350 5.475 1.755 ;
        RECT 9.885 1.350 10.055 1.755 ;
        RECT 14.465 1.350 14.635 1.755 ;
        RECT 19.045 1.350 19.215 1.755 ;
        RECT 0.490 1.050 21.750 1.350 ;
      LAYER mcon ;
        RECT 0.730 1.835 0.900 8.165 ;
        RECT 5.310 1.835 5.480 8.165 ;
        RECT 9.890 1.835 10.060 8.165 ;
        RECT 14.470 1.835 14.640 8.165 ;
        RECT 19.050 1.835 19.220 8.165 ;
      LAYER met1 ;
        RECT 0.700 1.775 0.930 8.225 ;
        RECT 5.280 1.775 5.510 8.225 ;
        RECT 9.860 1.775 10.090 8.225 ;
        RECT 14.440 1.775 14.670 8.225 ;
        RECT 19.020 1.775 19.250 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.470 21.750 9.700 ;
        RECT 0.490 1.465 21.750 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 21.750 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
        RECT 15.340 9.250 15.640 9.550 ;
        RECT 17.340 9.250 17.640 9.550 ;
        RECT 19.340 9.250 19.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 21.750 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 21.750 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
        RECT 15.340 -0.150 15.640 0.150 ;
        RECT 17.340 -0.150 17.640 0.150 ;
        RECT 19.340 -0.150 19.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 21.750 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9

#--------EOF---------

END LIBRARY