module macro (
    inout vdd,
    inout gnd,
    inout porst,
    inout va, 
    inout vb,
    inout vbg
 );
endmodule