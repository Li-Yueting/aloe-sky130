VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.800 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER met1 ;
        RECT 2.420 3.170 52.380 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 51.264000 ;
    PORT
      LAYER met1 ;
        RECT 1.550 6.750 53.250 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 107.630394 ;
    PORT
      LAYER pwell ;
        RECT 0.600 7.285 54.200 8.050 ;
        RECT 0.600 2.115 1.365 7.285 ;
        RECT 6.535 2.115 8.065 7.285 ;
        RECT 13.235 2.115 14.765 7.285 ;
        RECT 19.935 2.115 21.465 7.285 ;
        RECT 26.635 2.115 28.165 7.285 ;
        RECT 33.335 2.115 34.865 7.285 ;
        RECT 40.035 2.115 41.565 7.285 ;
        RECT 46.735 2.115 48.265 7.285 ;
        RECT 53.435 2.115 54.200 7.285 ;
        RECT 0.600 1.350 54.200 2.115 ;
      LAYER met1 ;
        RECT 0.730 7.500 54.070 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.600 9.100 54.200 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.600 -0.300 54.200 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.600 9.250 54.200 9.550 ;
        RECT 0.730 7.425 54.070 7.920 ;
        RECT 0.730 1.975 1.225 7.425 ;
        RECT 1.545 6.745 6.355 7.105 ;
        RECT 1.545 2.655 1.905 6.745 ;
        RECT 2.215 2.965 5.685 6.435 ;
        RECT 5.995 2.655 6.355 6.745 ;
        RECT 1.545 2.295 6.355 2.655 ;
        RECT 6.675 1.975 7.925 7.425 ;
        RECT 8.245 6.745 13.055 7.105 ;
        RECT 8.245 2.655 8.605 6.745 ;
        RECT 8.915 2.965 12.385 6.435 ;
        RECT 12.695 2.655 13.055 6.745 ;
        RECT 8.245 2.295 13.055 2.655 ;
        RECT 13.375 1.975 14.625 7.425 ;
        RECT 14.945 6.745 19.755 7.105 ;
        RECT 14.945 2.655 15.305 6.745 ;
        RECT 15.615 2.965 19.085 6.435 ;
        RECT 19.395 2.655 19.755 6.745 ;
        RECT 14.945 2.295 19.755 2.655 ;
        RECT 20.075 1.975 21.325 7.425 ;
        RECT 21.645 6.745 26.455 7.105 ;
        RECT 21.645 2.655 22.005 6.745 ;
        RECT 22.315 2.965 25.785 6.435 ;
        RECT 26.095 2.655 26.455 6.745 ;
        RECT 21.645 2.295 26.455 2.655 ;
        RECT 26.775 1.975 28.025 7.425 ;
        RECT 28.345 6.745 33.155 7.105 ;
        RECT 28.345 2.655 28.705 6.745 ;
        RECT 29.015 2.965 32.485 6.435 ;
        RECT 32.795 2.655 33.155 6.745 ;
        RECT 28.345 2.295 33.155 2.655 ;
        RECT 33.475 1.975 34.725 7.425 ;
        RECT 35.045 6.745 39.855 7.105 ;
        RECT 35.045 2.655 35.405 6.745 ;
        RECT 35.715 2.965 39.185 6.435 ;
        RECT 39.495 2.655 39.855 6.745 ;
        RECT 35.045 2.295 39.855 2.655 ;
        RECT 40.175 1.975 41.425 7.425 ;
        RECT 41.745 6.745 46.555 7.105 ;
        RECT 41.745 2.655 42.105 6.745 ;
        RECT 42.415 2.965 45.885 6.435 ;
        RECT 46.195 2.655 46.555 6.745 ;
        RECT 41.745 2.295 46.555 2.655 ;
        RECT 46.875 1.975 48.125 7.425 ;
        RECT 48.445 6.745 53.255 7.105 ;
        RECT 48.445 2.655 48.805 6.745 ;
        RECT 49.115 2.965 52.585 6.435 ;
        RECT 52.895 2.655 53.255 6.745 ;
        RECT 48.445 2.295 53.255 2.655 ;
        RECT 53.575 1.975 54.070 7.425 ;
        RECT 0.730 1.480 54.070 1.975 ;
        RECT 0.600 -0.150 54.200 0.150 ;
      LAYER mcon ;
        RECT 1.450 9.250 1.750 9.550 ;
        RECT 2.450 9.250 2.750 9.550 ;
        RECT 3.450 9.250 3.750 9.550 ;
        RECT 4.450 9.250 4.750 9.550 ;
        RECT 5.450 9.250 5.750 9.550 ;
        RECT 6.450 9.250 6.750 9.550 ;
        RECT 7.450 9.250 7.750 9.550 ;
        RECT 8.450 9.250 8.750 9.550 ;
        RECT 9.450 9.250 9.750 9.550 ;
        RECT 10.450 9.250 10.750 9.550 ;
        RECT 11.450 9.250 11.750 9.550 ;
        RECT 12.450 9.250 12.750 9.550 ;
        RECT 13.450 9.250 13.750 9.550 ;
        RECT 14.450 9.250 14.750 9.550 ;
        RECT 15.450 9.250 15.750 9.550 ;
        RECT 16.450 9.250 16.750 9.550 ;
        RECT 17.450 9.250 17.750 9.550 ;
        RECT 18.450 9.250 18.750 9.550 ;
        RECT 19.450 9.250 19.750 9.550 ;
        RECT 20.450 9.250 20.750 9.550 ;
        RECT 21.450 9.250 21.750 9.550 ;
        RECT 22.450 9.250 22.750 9.550 ;
        RECT 23.450 9.250 23.750 9.550 ;
        RECT 24.450 9.250 24.750 9.550 ;
        RECT 25.450 9.250 25.750 9.550 ;
        RECT 26.450 9.250 26.750 9.550 ;
        RECT 27.450 9.250 27.750 9.550 ;
        RECT 28.450 9.250 28.750 9.550 ;
        RECT 29.450 9.250 29.750 9.550 ;
        RECT 30.450 9.250 30.750 9.550 ;
        RECT 31.450 9.250 31.750 9.550 ;
        RECT 32.450 9.250 32.750 9.550 ;
        RECT 33.450 9.250 33.750 9.550 ;
        RECT 34.450 9.250 34.750 9.550 ;
        RECT 35.450 9.250 35.750 9.550 ;
        RECT 36.450 9.250 36.750 9.550 ;
        RECT 37.450 9.250 37.750 9.550 ;
        RECT 38.450 9.250 38.750 9.550 ;
        RECT 39.450 9.250 39.750 9.550 ;
        RECT 40.450 9.250 40.750 9.550 ;
        RECT 41.450 9.250 41.750 9.550 ;
        RECT 42.450 9.250 42.750 9.550 ;
        RECT 43.450 9.250 43.750 9.550 ;
        RECT 44.450 9.250 44.750 9.550 ;
        RECT 45.450 9.250 45.750 9.550 ;
        RECT 46.450 9.250 46.750 9.550 ;
        RECT 47.450 9.250 47.750 9.550 ;
        RECT 48.450 9.250 48.750 9.550 ;
        RECT 49.450 9.250 49.750 9.550 ;
        RECT 50.450 9.250 50.750 9.550 ;
        RECT 51.450 9.250 51.750 9.550 ;
        RECT 52.450 9.250 52.750 9.550 ;
        RECT 53.450 9.250 53.750 9.550 ;
        RECT 0.830 7.650 1.000 7.820 ;
        RECT 1.280 7.650 1.450 7.820 ;
        RECT 1.730 7.650 1.900 7.820 ;
        RECT 2.180 7.650 2.350 7.820 ;
        RECT 2.630 7.650 2.800 7.820 ;
        RECT 3.080 7.650 3.250 7.820 ;
        RECT 3.530 7.650 3.700 7.820 ;
        RECT 3.980 7.650 4.150 7.820 ;
        RECT 4.430 7.650 4.600 7.820 ;
        RECT 4.880 7.650 5.050 7.820 ;
        RECT 5.330 7.650 5.500 7.820 ;
        RECT 5.780 7.650 5.950 7.820 ;
        RECT 6.230 7.650 6.400 7.820 ;
        RECT 6.680 7.650 6.850 7.820 ;
        RECT 7.530 7.650 7.700 7.820 ;
        RECT 7.980 7.650 8.150 7.820 ;
        RECT 8.430 7.650 8.600 7.820 ;
        RECT 8.880 7.650 9.050 7.820 ;
        RECT 9.330 7.650 9.500 7.820 ;
        RECT 9.780 7.650 9.950 7.820 ;
        RECT 10.230 7.650 10.400 7.820 ;
        RECT 10.680 7.650 10.850 7.820 ;
        RECT 11.130 7.650 11.300 7.820 ;
        RECT 11.580 7.650 11.750 7.820 ;
        RECT 12.030 7.650 12.200 7.820 ;
        RECT 12.480 7.650 12.650 7.820 ;
        RECT 12.930 7.650 13.100 7.820 ;
        RECT 13.380 7.650 13.550 7.820 ;
        RECT 14.230 7.650 14.400 7.820 ;
        RECT 14.680 7.650 14.850 7.820 ;
        RECT 15.130 7.650 15.300 7.820 ;
        RECT 15.580 7.650 15.750 7.820 ;
        RECT 16.030 7.650 16.200 7.820 ;
        RECT 16.480 7.650 16.650 7.820 ;
        RECT 16.930 7.650 17.100 7.820 ;
        RECT 17.380 7.650 17.550 7.820 ;
        RECT 17.830 7.650 18.000 7.820 ;
        RECT 18.280 7.650 18.450 7.820 ;
        RECT 18.730 7.650 18.900 7.820 ;
        RECT 19.180 7.650 19.350 7.820 ;
        RECT 19.630 7.650 19.800 7.820 ;
        RECT 20.080 7.650 20.250 7.820 ;
        RECT 20.930 7.650 21.100 7.820 ;
        RECT 21.380 7.650 21.550 7.820 ;
        RECT 21.830 7.650 22.000 7.820 ;
        RECT 22.280 7.650 22.450 7.820 ;
        RECT 22.730 7.650 22.900 7.820 ;
        RECT 23.180 7.650 23.350 7.820 ;
        RECT 23.630 7.650 23.800 7.820 ;
        RECT 24.080 7.650 24.250 7.820 ;
        RECT 24.530 7.650 24.700 7.820 ;
        RECT 24.980 7.650 25.150 7.820 ;
        RECT 25.430 7.650 25.600 7.820 ;
        RECT 25.880 7.650 26.050 7.820 ;
        RECT 26.330 7.650 26.500 7.820 ;
        RECT 26.780 7.650 26.950 7.820 ;
        RECT 27.630 7.650 27.800 7.820 ;
        RECT 28.080 7.650 28.250 7.820 ;
        RECT 28.530 7.650 28.700 7.820 ;
        RECT 28.980 7.650 29.150 7.820 ;
        RECT 29.430 7.650 29.600 7.820 ;
        RECT 29.880 7.650 30.050 7.820 ;
        RECT 30.330 7.650 30.500 7.820 ;
        RECT 30.780 7.650 30.950 7.820 ;
        RECT 31.230 7.650 31.400 7.820 ;
        RECT 31.680 7.650 31.850 7.820 ;
        RECT 32.130 7.650 32.300 7.820 ;
        RECT 32.580 7.650 32.750 7.820 ;
        RECT 33.030 7.650 33.200 7.820 ;
        RECT 33.480 7.650 33.650 7.820 ;
        RECT 34.330 7.650 34.500 7.820 ;
        RECT 34.780 7.650 34.950 7.820 ;
        RECT 35.230 7.650 35.400 7.820 ;
        RECT 35.680 7.650 35.850 7.820 ;
        RECT 36.130 7.650 36.300 7.820 ;
        RECT 36.580 7.650 36.750 7.820 ;
        RECT 37.030 7.650 37.200 7.820 ;
        RECT 37.480 7.650 37.650 7.820 ;
        RECT 37.930 7.650 38.100 7.820 ;
        RECT 38.380 7.650 38.550 7.820 ;
        RECT 38.830 7.650 39.000 7.820 ;
        RECT 39.280 7.650 39.450 7.820 ;
        RECT 39.730 7.650 39.900 7.820 ;
        RECT 40.180 7.650 40.350 7.820 ;
        RECT 41.030 7.650 41.200 7.820 ;
        RECT 41.480 7.650 41.650 7.820 ;
        RECT 41.930 7.650 42.100 7.820 ;
        RECT 42.380 7.650 42.550 7.820 ;
        RECT 42.830 7.650 43.000 7.820 ;
        RECT 43.280 7.650 43.450 7.820 ;
        RECT 43.730 7.650 43.900 7.820 ;
        RECT 44.180 7.650 44.350 7.820 ;
        RECT 44.630 7.650 44.800 7.820 ;
        RECT 45.080 7.650 45.250 7.820 ;
        RECT 45.530 7.650 45.700 7.820 ;
        RECT 45.980 7.650 46.150 7.820 ;
        RECT 46.430 7.650 46.600 7.820 ;
        RECT 46.880 7.650 47.050 7.820 ;
        RECT 47.730 7.650 47.900 7.820 ;
        RECT 48.180 7.650 48.350 7.820 ;
        RECT 48.630 7.650 48.800 7.820 ;
        RECT 49.080 7.650 49.250 7.820 ;
        RECT 49.530 7.650 49.700 7.820 ;
        RECT 49.980 7.650 50.150 7.820 ;
        RECT 50.430 7.650 50.600 7.820 ;
        RECT 50.880 7.650 51.050 7.820 ;
        RECT 51.330 7.650 51.500 7.820 ;
        RECT 51.780 7.650 51.950 7.820 ;
        RECT 52.230 7.650 52.400 7.820 ;
        RECT 52.680 7.650 52.850 7.820 ;
        RECT 53.130 7.650 53.300 7.820 ;
        RECT 53.580 7.650 53.750 7.820 ;
        RECT 1.650 6.850 1.820 7.020 ;
        RECT 2.100 6.850 2.270 7.020 ;
        RECT 2.550 6.850 2.720 7.020 ;
        RECT 3.000 6.850 3.170 7.020 ;
        RECT 3.450 6.850 3.620 7.020 ;
        RECT 3.900 6.850 4.070 7.020 ;
        RECT 4.350 6.850 4.520 7.020 ;
        RECT 4.800 6.850 4.970 7.020 ;
        RECT 5.250 6.850 5.420 7.020 ;
        RECT 5.700 6.850 5.870 7.020 ;
        RECT 6.150 6.850 6.320 7.020 ;
        RECT 2.580 5.830 2.750 6.000 ;
        RECT 3.080 5.830 3.250 6.000 ;
        RECT 3.580 5.830 3.750 6.000 ;
        RECT 4.080 5.830 4.250 6.000 ;
        RECT 4.580 5.830 4.750 6.000 ;
        RECT 5.080 5.830 5.250 6.000 ;
        RECT 2.580 5.330 2.750 5.500 ;
        RECT 3.080 5.330 3.250 5.500 ;
        RECT 3.580 5.330 3.750 5.500 ;
        RECT 4.080 5.330 4.250 5.500 ;
        RECT 4.580 5.330 4.750 5.500 ;
        RECT 5.080 5.330 5.250 5.500 ;
        RECT 2.580 4.830 2.750 5.000 ;
        RECT 3.080 4.830 3.250 5.000 ;
        RECT 3.580 4.830 3.750 5.000 ;
        RECT 4.080 4.830 4.250 5.000 ;
        RECT 4.580 4.830 4.750 5.000 ;
        RECT 5.080 4.830 5.250 5.000 ;
        RECT 2.580 4.330 2.750 4.500 ;
        RECT 3.080 4.330 3.250 4.500 ;
        RECT 3.580 4.330 3.750 4.500 ;
        RECT 4.080 4.330 4.250 4.500 ;
        RECT 4.580 4.330 4.750 4.500 ;
        RECT 5.080 4.330 5.250 4.500 ;
        RECT 2.580 3.830 2.750 4.000 ;
        RECT 3.080 3.830 3.250 4.000 ;
        RECT 3.580 3.830 3.750 4.000 ;
        RECT 4.080 3.830 4.250 4.000 ;
        RECT 4.580 3.830 4.750 4.000 ;
        RECT 5.080 3.830 5.250 4.000 ;
        RECT 2.580 3.330 2.750 3.500 ;
        RECT 3.080 3.330 3.250 3.500 ;
        RECT 3.580 3.330 3.750 3.500 ;
        RECT 4.080 3.330 4.250 3.500 ;
        RECT 4.580 3.330 4.750 3.500 ;
        RECT 5.080 3.330 5.250 3.500 ;
        RECT 8.350 6.850 8.520 7.020 ;
        RECT 8.800 6.850 8.970 7.020 ;
        RECT 9.250 6.850 9.420 7.020 ;
        RECT 9.700 6.850 9.870 7.020 ;
        RECT 10.150 6.850 10.320 7.020 ;
        RECT 10.600 6.850 10.770 7.020 ;
        RECT 11.050 6.850 11.220 7.020 ;
        RECT 11.500 6.850 11.670 7.020 ;
        RECT 11.950 6.850 12.120 7.020 ;
        RECT 12.400 6.850 12.570 7.020 ;
        RECT 12.850 6.850 13.020 7.020 ;
        RECT 9.280 5.830 9.450 6.000 ;
        RECT 9.780 5.830 9.950 6.000 ;
        RECT 10.280 5.830 10.450 6.000 ;
        RECT 10.780 5.830 10.950 6.000 ;
        RECT 11.280 5.830 11.450 6.000 ;
        RECT 11.780 5.830 11.950 6.000 ;
        RECT 9.280 5.330 9.450 5.500 ;
        RECT 9.780 5.330 9.950 5.500 ;
        RECT 10.280 5.330 10.450 5.500 ;
        RECT 10.780 5.330 10.950 5.500 ;
        RECT 11.280 5.330 11.450 5.500 ;
        RECT 11.780 5.330 11.950 5.500 ;
        RECT 9.280 4.830 9.450 5.000 ;
        RECT 9.780 4.830 9.950 5.000 ;
        RECT 10.280 4.830 10.450 5.000 ;
        RECT 10.780 4.830 10.950 5.000 ;
        RECT 11.280 4.830 11.450 5.000 ;
        RECT 11.780 4.830 11.950 5.000 ;
        RECT 9.280 4.330 9.450 4.500 ;
        RECT 9.780 4.330 9.950 4.500 ;
        RECT 10.280 4.330 10.450 4.500 ;
        RECT 10.780 4.330 10.950 4.500 ;
        RECT 11.280 4.330 11.450 4.500 ;
        RECT 11.780 4.330 11.950 4.500 ;
        RECT 9.280 3.830 9.450 4.000 ;
        RECT 9.780 3.830 9.950 4.000 ;
        RECT 10.280 3.830 10.450 4.000 ;
        RECT 10.780 3.830 10.950 4.000 ;
        RECT 11.280 3.830 11.450 4.000 ;
        RECT 11.780 3.830 11.950 4.000 ;
        RECT 9.280 3.330 9.450 3.500 ;
        RECT 9.780 3.330 9.950 3.500 ;
        RECT 10.280 3.330 10.450 3.500 ;
        RECT 10.780 3.330 10.950 3.500 ;
        RECT 11.280 3.330 11.450 3.500 ;
        RECT 11.780 3.330 11.950 3.500 ;
        RECT 15.050 6.850 15.220 7.020 ;
        RECT 15.500 6.850 15.670 7.020 ;
        RECT 15.950 6.850 16.120 7.020 ;
        RECT 16.400 6.850 16.570 7.020 ;
        RECT 16.850 6.850 17.020 7.020 ;
        RECT 17.300 6.850 17.470 7.020 ;
        RECT 17.750 6.850 17.920 7.020 ;
        RECT 18.200 6.850 18.370 7.020 ;
        RECT 18.650 6.850 18.820 7.020 ;
        RECT 19.100 6.850 19.270 7.020 ;
        RECT 19.550 6.850 19.720 7.020 ;
        RECT 15.980 5.830 16.150 6.000 ;
        RECT 16.480 5.830 16.650 6.000 ;
        RECT 16.980 5.830 17.150 6.000 ;
        RECT 17.480 5.830 17.650 6.000 ;
        RECT 17.980 5.830 18.150 6.000 ;
        RECT 18.480 5.830 18.650 6.000 ;
        RECT 15.980 5.330 16.150 5.500 ;
        RECT 16.480 5.330 16.650 5.500 ;
        RECT 16.980 5.330 17.150 5.500 ;
        RECT 17.480 5.330 17.650 5.500 ;
        RECT 17.980 5.330 18.150 5.500 ;
        RECT 18.480 5.330 18.650 5.500 ;
        RECT 15.980 4.830 16.150 5.000 ;
        RECT 16.480 4.830 16.650 5.000 ;
        RECT 16.980 4.830 17.150 5.000 ;
        RECT 17.480 4.830 17.650 5.000 ;
        RECT 17.980 4.830 18.150 5.000 ;
        RECT 18.480 4.830 18.650 5.000 ;
        RECT 15.980 4.330 16.150 4.500 ;
        RECT 16.480 4.330 16.650 4.500 ;
        RECT 16.980 4.330 17.150 4.500 ;
        RECT 17.480 4.330 17.650 4.500 ;
        RECT 17.980 4.330 18.150 4.500 ;
        RECT 18.480 4.330 18.650 4.500 ;
        RECT 15.980 3.830 16.150 4.000 ;
        RECT 16.480 3.830 16.650 4.000 ;
        RECT 16.980 3.830 17.150 4.000 ;
        RECT 17.480 3.830 17.650 4.000 ;
        RECT 17.980 3.830 18.150 4.000 ;
        RECT 18.480 3.830 18.650 4.000 ;
        RECT 15.980 3.330 16.150 3.500 ;
        RECT 16.480 3.330 16.650 3.500 ;
        RECT 16.980 3.330 17.150 3.500 ;
        RECT 17.480 3.330 17.650 3.500 ;
        RECT 17.980 3.330 18.150 3.500 ;
        RECT 18.480 3.330 18.650 3.500 ;
        RECT 21.750 6.850 21.920 7.020 ;
        RECT 22.200 6.850 22.370 7.020 ;
        RECT 22.650 6.850 22.820 7.020 ;
        RECT 23.100 6.850 23.270 7.020 ;
        RECT 23.550 6.850 23.720 7.020 ;
        RECT 24.000 6.850 24.170 7.020 ;
        RECT 24.450 6.850 24.620 7.020 ;
        RECT 24.900 6.850 25.070 7.020 ;
        RECT 25.350 6.850 25.520 7.020 ;
        RECT 25.800 6.850 25.970 7.020 ;
        RECT 26.250 6.850 26.420 7.020 ;
        RECT 22.680 5.830 22.850 6.000 ;
        RECT 23.180 5.830 23.350 6.000 ;
        RECT 23.680 5.830 23.850 6.000 ;
        RECT 24.180 5.830 24.350 6.000 ;
        RECT 24.680 5.830 24.850 6.000 ;
        RECT 25.180 5.830 25.350 6.000 ;
        RECT 22.680 5.330 22.850 5.500 ;
        RECT 23.180 5.330 23.350 5.500 ;
        RECT 23.680 5.330 23.850 5.500 ;
        RECT 24.180 5.330 24.350 5.500 ;
        RECT 24.680 5.330 24.850 5.500 ;
        RECT 25.180 5.330 25.350 5.500 ;
        RECT 22.680 4.830 22.850 5.000 ;
        RECT 23.180 4.830 23.350 5.000 ;
        RECT 23.680 4.830 23.850 5.000 ;
        RECT 24.180 4.830 24.350 5.000 ;
        RECT 24.680 4.830 24.850 5.000 ;
        RECT 25.180 4.830 25.350 5.000 ;
        RECT 22.680 4.330 22.850 4.500 ;
        RECT 23.180 4.330 23.350 4.500 ;
        RECT 23.680 4.330 23.850 4.500 ;
        RECT 24.180 4.330 24.350 4.500 ;
        RECT 24.680 4.330 24.850 4.500 ;
        RECT 25.180 4.330 25.350 4.500 ;
        RECT 22.680 3.830 22.850 4.000 ;
        RECT 23.180 3.830 23.350 4.000 ;
        RECT 23.680 3.830 23.850 4.000 ;
        RECT 24.180 3.830 24.350 4.000 ;
        RECT 24.680 3.830 24.850 4.000 ;
        RECT 25.180 3.830 25.350 4.000 ;
        RECT 22.680 3.330 22.850 3.500 ;
        RECT 23.180 3.330 23.350 3.500 ;
        RECT 23.680 3.330 23.850 3.500 ;
        RECT 24.180 3.330 24.350 3.500 ;
        RECT 24.680 3.330 24.850 3.500 ;
        RECT 25.180 3.330 25.350 3.500 ;
        RECT 28.450 6.850 28.620 7.020 ;
        RECT 28.900 6.850 29.070 7.020 ;
        RECT 29.350 6.850 29.520 7.020 ;
        RECT 29.800 6.850 29.970 7.020 ;
        RECT 30.250 6.850 30.420 7.020 ;
        RECT 30.700 6.850 30.870 7.020 ;
        RECT 31.150 6.850 31.320 7.020 ;
        RECT 31.600 6.850 31.770 7.020 ;
        RECT 32.050 6.850 32.220 7.020 ;
        RECT 32.500 6.850 32.670 7.020 ;
        RECT 32.950 6.850 33.120 7.020 ;
        RECT 29.380 5.830 29.550 6.000 ;
        RECT 29.880 5.830 30.050 6.000 ;
        RECT 30.380 5.830 30.550 6.000 ;
        RECT 30.880 5.830 31.050 6.000 ;
        RECT 31.380 5.830 31.550 6.000 ;
        RECT 31.880 5.830 32.050 6.000 ;
        RECT 29.380 5.330 29.550 5.500 ;
        RECT 29.880 5.330 30.050 5.500 ;
        RECT 30.380 5.330 30.550 5.500 ;
        RECT 30.880 5.330 31.050 5.500 ;
        RECT 31.380 5.330 31.550 5.500 ;
        RECT 31.880 5.330 32.050 5.500 ;
        RECT 29.380 4.830 29.550 5.000 ;
        RECT 29.880 4.830 30.050 5.000 ;
        RECT 30.380 4.830 30.550 5.000 ;
        RECT 30.880 4.830 31.050 5.000 ;
        RECT 31.380 4.830 31.550 5.000 ;
        RECT 31.880 4.830 32.050 5.000 ;
        RECT 29.380 4.330 29.550 4.500 ;
        RECT 29.880 4.330 30.050 4.500 ;
        RECT 30.380 4.330 30.550 4.500 ;
        RECT 30.880 4.330 31.050 4.500 ;
        RECT 31.380 4.330 31.550 4.500 ;
        RECT 31.880 4.330 32.050 4.500 ;
        RECT 29.380 3.830 29.550 4.000 ;
        RECT 29.880 3.830 30.050 4.000 ;
        RECT 30.380 3.830 30.550 4.000 ;
        RECT 30.880 3.830 31.050 4.000 ;
        RECT 31.380 3.830 31.550 4.000 ;
        RECT 31.880 3.830 32.050 4.000 ;
        RECT 29.380 3.330 29.550 3.500 ;
        RECT 29.880 3.330 30.050 3.500 ;
        RECT 30.380 3.330 30.550 3.500 ;
        RECT 30.880 3.330 31.050 3.500 ;
        RECT 31.380 3.330 31.550 3.500 ;
        RECT 31.880 3.330 32.050 3.500 ;
        RECT 35.150 6.850 35.320 7.020 ;
        RECT 35.600 6.850 35.770 7.020 ;
        RECT 36.050 6.850 36.220 7.020 ;
        RECT 36.500 6.850 36.670 7.020 ;
        RECT 36.950 6.850 37.120 7.020 ;
        RECT 37.400 6.850 37.570 7.020 ;
        RECT 37.850 6.850 38.020 7.020 ;
        RECT 38.300 6.850 38.470 7.020 ;
        RECT 38.750 6.850 38.920 7.020 ;
        RECT 39.200 6.850 39.370 7.020 ;
        RECT 39.650 6.850 39.820 7.020 ;
        RECT 36.080 5.830 36.250 6.000 ;
        RECT 36.580 5.830 36.750 6.000 ;
        RECT 37.080 5.830 37.250 6.000 ;
        RECT 37.580 5.830 37.750 6.000 ;
        RECT 38.080 5.830 38.250 6.000 ;
        RECT 38.580 5.830 38.750 6.000 ;
        RECT 36.080 5.330 36.250 5.500 ;
        RECT 36.580 5.330 36.750 5.500 ;
        RECT 37.080 5.330 37.250 5.500 ;
        RECT 37.580 5.330 37.750 5.500 ;
        RECT 38.080 5.330 38.250 5.500 ;
        RECT 38.580 5.330 38.750 5.500 ;
        RECT 36.080 4.830 36.250 5.000 ;
        RECT 36.580 4.830 36.750 5.000 ;
        RECT 37.080 4.830 37.250 5.000 ;
        RECT 37.580 4.830 37.750 5.000 ;
        RECT 38.080 4.830 38.250 5.000 ;
        RECT 38.580 4.830 38.750 5.000 ;
        RECT 36.080 4.330 36.250 4.500 ;
        RECT 36.580 4.330 36.750 4.500 ;
        RECT 37.080 4.330 37.250 4.500 ;
        RECT 37.580 4.330 37.750 4.500 ;
        RECT 38.080 4.330 38.250 4.500 ;
        RECT 38.580 4.330 38.750 4.500 ;
        RECT 36.080 3.830 36.250 4.000 ;
        RECT 36.580 3.830 36.750 4.000 ;
        RECT 37.080 3.830 37.250 4.000 ;
        RECT 37.580 3.830 37.750 4.000 ;
        RECT 38.080 3.830 38.250 4.000 ;
        RECT 38.580 3.830 38.750 4.000 ;
        RECT 36.080 3.330 36.250 3.500 ;
        RECT 36.580 3.330 36.750 3.500 ;
        RECT 37.080 3.330 37.250 3.500 ;
        RECT 37.580 3.330 37.750 3.500 ;
        RECT 38.080 3.330 38.250 3.500 ;
        RECT 38.580 3.330 38.750 3.500 ;
        RECT 41.850 6.850 42.020 7.020 ;
        RECT 42.300 6.850 42.470 7.020 ;
        RECT 42.750 6.850 42.920 7.020 ;
        RECT 43.200 6.850 43.370 7.020 ;
        RECT 43.650 6.850 43.820 7.020 ;
        RECT 44.100 6.850 44.270 7.020 ;
        RECT 44.550 6.850 44.720 7.020 ;
        RECT 45.000 6.850 45.170 7.020 ;
        RECT 45.450 6.850 45.620 7.020 ;
        RECT 45.900 6.850 46.070 7.020 ;
        RECT 46.350 6.850 46.520 7.020 ;
        RECT 42.780 5.830 42.950 6.000 ;
        RECT 43.280 5.830 43.450 6.000 ;
        RECT 43.780 5.830 43.950 6.000 ;
        RECT 44.280 5.830 44.450 6.000 ;
        RECT 44.780 5.830 44.950 6.000 ;
        RECT 45.280 5.830 45.450 6.000 ;
        RECT 42.780 5.330 42.950 5.500 ;
        RECT 43.280 5.330 43.450 5.500 ;
        RECT 43.780 5.330 43.950 5.500 ;
        RECT 44.280 5.330 44.450 5.500 ;
        RECT 44.780 5.330 44.950 5.500 ;
        RECT 45.280 5.330 45.450 5.500 ;
        RECT 42.780 4.830 42.950 5.000 ;
        RECT 43.280 4.830 43.450 5.000 ;
        RECT 43.780 4.830 43.950 5.000 ;
        RECT 44.280 4.830 44.450 5.000 ;
        RECT 44.780 4.830 44.950 5.000 ;
        RECT 45.280 4.830 45.450 5.000 ;
        RECT 42.780 4.330 42.950 4.500 ;
        RECT 43.280 4.330 43.450 4.500 ;
        RECT 43.780 4.330 43.950 4.500 ;
        RECT 44.280 4.330 44.450 4.500 ;
        RECT 44.780 4.330 44.950 4.500 ;
        RECT 45.280 4.330 45.450 4.500 ;
        RECT 42.780 3.830 42.950 4.000 ;
        RECT 43.280 3.830 43.450 4.000 ;
        RECT 43.780 3.830 43.950 4.000 ;
        RECT 44.280 3.830 44.450 4.000 ;
        RECT 44.780 3.830 44.950 4.000 ;
        RECT 45.280 3.830 45.450 4.000 ;
        RECT 42.780 3.330 42.950 3.500 ;
        RECT 43.280 3.330 43.450 3.500 ;
        RECT 43.780 3.330 43.950 3.500 ;
        RECT 44.280 3.330 44.450 3.500 ;
        RECT 44.780 3.330 44.950 3.500 ;
        RECT 45.280 3.330 45.450 3.500 ;
        RECT 48.550 6.850 48.720 7.020 ;
        RECT 49.000 6.850 49.170 7.020 ;
        RECT 49.450 6.850 49.620 7.020 ;
        RECT 49.900 6.850 50.070 7.020 ;
        RECT 50.350 6.850 50.520 7.020 ;
        RECT 50.800 6.850 50.970 7.020 ;
        RECT 51.250 6.850 51.420 7.020 ;
        RECT 51.700 6.850 51.870 7.020 ;
        RECT 52.150 6.850 52.320 7.020 ;
        RECT 52.600 6.850 52.770 7.020 ;
        RECT 53.050 6.850 53.220 7.020 ;
        RECT 49.480 5.830 49.650 6.000 ;
        RECT 49.980 5.830 50.150 6.000 ;
        RECT 50.480 5.830 50.650 6.000 ;
        RECT 50.980 5.830 51.150 6.000 ;
        RECT 51.480 5.830 51.650 6.000 ;
        RECT 51.980 5.830 52.150 6.000 ;
        RECT 49.480 5.330 49.650 5.500 ;
        RECT 49.980 5.330 50.150 5.500 ;
        RECT 50.480 5.330 50.650 5.500 ;
        RECT 50.980 5.330 51.150 5.500 ;
        RECT 51.480 5.330 51.650 5.500 ;
        RECT 51.980 5.330 52.150 5.500 ;
        RECT 49.480 4.830 49.650 5.000 ;
        RECT 49.980 4.830 50.150 5.000 ;
        RECT 50.480 4.830 50.650 5.000 ;
        RECT 50.980 4.830 51.150 5.000 ;
        RECT 51.480 4.830 51.650 5.000 ;
        RECT 51.980 4.830 52.150 5.000 ;
        RECT 49.480 4.330 49.650 4.500 ;
        RECT 49.980 4.330 50.150 4.500 ;
        RECT 50.480 4.330 50.650 4.500 ;
        RECT 50.980 4.330 51.150 4.500 ;
        RECT 51.480 4.330 51.650 4.500 ;
        RECT 51.980 4.330 52.150 4.500 ;
        RECT 49.480 3.830 49.650 4.000 ;
        RECT 49.980 3.830 50.150 4.000 ;
        RECT 50.480 3.830 50.650 4.000 ;
        RECT 50.980 3.830 51.150 4.000 ;
        RECT 51.480 3.830 51.650 4.000 ;
        RECT 51.980 3.830 52.150 4.000 ;
        RECT 49.480 3.330 49.650 3.500 ;
        RECT 49.980 3.330 50.150 3.500 ;
        RECT 50.480 3.330 50.650 3.500 ;
        RECT 50.980 3.330 51.150 3.500 ;
        RECT 51.480 3.330 51.650 3.500 ;
        RECT 51.980 3.330 52.150 3.500 ;
        RECT 1.450 -0.150 1.750 0.150 ;
        RECT 2.450 -0.150 2.750 0.150 ;
        RECT 3.450 -0.150 3.750 0.150 ;
        RECT 4.450 -0.150 4.750 0.150 ;
        RECT 5.450 -0.150 5.750 0.150 ;
        RECT 6.450 -0.150 6.750 0.150 ;
        RECT 7.450 -0.150 7.750 0.150 ;
        RECT 8.450 -0.150 8.750 0.150 ;
        RECT 9.450 -0.150 9.750 0.150 ;
        RECT 10.450 -0.150 10.750 0.150 ;
        RECT 11.450 -0.150 11.750 0.150 ;
        RECT 12.450 -0.150 12.750 0.150 ;
        RECT 13.450 -0.150 13.750 0.150 ;
        RECT 14.450 -0.150 14.750 0.150 ;
        RECT 15.450 -0.150 15.750 0.150 ;
        RECT 16.450 -0.150 16.750 0.150 ;
        RECT 17.450 -0.150 17.750 0.150 ;
        RECT 18.450 -0.150 18.750 0.150 ;
        RECT 19.450 -0.150 19.750 0.150 ;
        RECT 20.450 -0.150 20.750 0.150 ;
        RECT 21.450 -0.150 21.750 0.150 ;
        RECT 22.450 -0.150 22.750 0.150 ;
        RECT 23.450 -0.150 23.750 0.150 ;
        RECT 24.450 -0.150 24.750 0.150 ;
        RECT 25.450 -0.150 25.750 0.150 ;
        RECT 26.450 -0.150 26.750 0.150 ;
        RECT 27.450 -0.150 27.750 0.150 ;
        RECT 28.450 -0.150 28.750 0.150 ;
        RECT 29.450 -0.150 29.750 0.150 ;
        RECT 30.450 -0.150 30.750 0.150 ;
        RECT 31.450 -0.150 31.750 0.150 ;
        RECT 32.450 -0.150 32.750 0.150 ;
        RECT 33.450 -0.150 33.750 0.150 ;
        RECT 34.450 -0.150 34.750 0.150 ;
        RECT 35.450 -0.150 35.750 0.150 ;
        RECT 36.450 -0.150 36.750 0.150 ;
        RECT 37.450 -0.150 37.750 0.150 ;
        RECT 38.450 -0.150 38.750 0.150 ;
        RECT 39.450 -0.150 39.750 0.150 ;
        RECT 40.450 -0.150 40.750 0.150 ;
        RECT 41.450 -0.150 41.750 0.150 ;
        RECT 42.450 -0.150 42.750 0.150 ;
        RECT 43.450 -0.150 43.750 0.150 ;
        RECT 44.450 -0.150 44.750 0.150 ;
        RECT 45.450 -0.150 45.750 0.150 ;
        RECT 46.450 -0.150 46.750 0.150 ;
        RECT 47.450 -0.150 47.750 0.150 ;
        RECT 48.450 -0.150 48.750 0.150 ;
        RECT 49.450 -0.150 49.750 0.150 ;
        RECT 50.450 -0.150 50.750 0.150 ;
        RECT 51.450 -0.150 51.750 0.150 ;
        RECT 52.450 -0.150 52.750 0.150 ;
        RECT 53.450 -0.150 53.750 0.150 ;
  END
END sky130_asc_pnp_05v5_W3p40L3p40_8

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.970 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.340 0.720 3.520 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 8.450 3.520 8.750 ;
        RECT 3.285 7.020 3.455 8.450 ;
        RECT 3.285 6.930 3.460 7.020 ;
        RECT 3.290 2.980 3.460 6.930 ;
      LAYER mcon ;
        RECT 3.290 3.060 3.460 6.940 ;
      LAYER met1 ;
        RECT 3.260 3.000 3.490 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 1.000 3.270 1.170 7.020 ;
        RECT 0.995 2.980 1.170 3.270 ;
        RECT 0.995 2.150 1.165 2.980 ;
        RECT 0.940 1.850 3.520 2.150 ;
      LAYER mcon ;
        RECT 1.000 3.060 1.170 6.940 ;
      LAYER met1 ;
        RECT 0.970 3.000 1.200 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 3.520 9.550 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 3.520 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.450 0.150 3.520 7.130 ;
      LAYER li1 ;
        RECT 0.590 0.150 0.890 1.200 ;
        RECT 0.450 -0.150 3.520 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 3.520 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.630 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 4.030 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 4.030 8.650 ;
        RECT 3.615 8.245 3.785 8.450 ;
        RECT 3.615 8.130 3.790 8.245 ;
        RECT 3.620 1.755 3.790 8.130 ;
      LAYER mcon ;
        RECT 3.620 1.835 3.790 8.165 ;
      LAYER met1 ;
        RECT 3.590 1.775 3.820 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 1.330 1.870 1.500 8.245 ;
        RECT 1.325 1.755 1.500 1.870 ;
        RECT 1.325 1.350 1.495 1.755 ;
        RECT 1.090 1.050 4.030 1.350 ;
      LAYER mcon ;
        RECT 1.330 1.835 1.500 8.165 ;
      LAYER met1 ;
        RECT 1.300 1.775 1.530 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 1.470 4.030 9.700 ;
        RECT 1.090 1.465 4.030 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 4.030 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 4.030 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 4.030 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 4.030 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_res_xhigh_po_2p85_1
  CLASS CORE ;
  FOREIGN sky130_asc_res_xhigh_po_2p85_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.600 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 0.755 5.395 2.805 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 0.755 0.595 2.805 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.700 9.100 12.900 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.700 -0.300 12.900 8.250 ;
      LAYER met1 ;
        RECT 0.700 -0.300 12.900 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.700 9.250 12.900 9.550 ;
        RECT 0.700 5.375 2.860 8.225 ;
        RECT 0.700 0.575 2.860 3.425 ;
        RECT 5.260 0.150 8.340 4.850 ;
        RECT 10.740 0.575 12.900 8.225 ;
        RECT 0.700 -0.150 12.900 0.150 ;
      LAYER mcon ;
        RECT 1.550 9.250 1.850 9.550 ;
        RECT 2.550 9.250 2.850 9.550 ;
        RECT 3.550 9.250 3.850 9.550 ;
        RECT 4.550 9.250 4.850 9.550 ;
        RECT 5.550 9.250 5.850 9.550 ;
        RECT 6.550 9.250 6.850 9.550 ;
        RECT 7.550 9.250 7.850 9.550 ;
        RECT 8.550 9.250 8.850 9.550 ;
        RECT 9.550 9.250 9.850 9.550 ;
        RECT 10.550 9.250 10.850 9.550 ;
        RECT 11.550 9.250 11.850 9.550 ;
        RECT 0.790 5.455 2.775 8.145 ;
        RECT 10.825 5.455 12.810 8.145 ;
        RECT 0.790 0.655 2.775 3.345 ;
        RECT 10.825 0.655 12.810 3.345 ;
        RECT 1.550 -0.150 1.850 0.150 ;
        RECT 2.550 -0.150 2.850 0.150 ;
        RECT 3.550 -0.150 3.850 0.150 ;
        RECT 4.550 -0.150 4.850 0.150 ;
        RECT 5.550 -0.150 5.850 0.150 ;
        RECT 6.550 -0.150 6.850 0.150 ;
        RECT 7.550 -0.150 7.850 0.150 ;
        RECT 8.550 -0.150 8.850 0.150 ;
        RECT 9.550 -0.150 9.850 0.150 ;
        RECT 10.550 -0.150 10.850 0.150 ;
        RECT 11.550 -0.150 11.850 0.150 ;
      LAYER met1 ;
        RECT 10.795 5.395 12.845 8.205 ;
        RECT 10.740 0.575 12.900 5.395 ;
  END
END sky130_asc_res_xhigh_po_2p85_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 139.735 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 139.130 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 139.130 8.650 ;
        RECT 3.615 1.755 3.785 8.450 ;
        RECT 8.195 1.755 8.365 8.450 ;
        RECT 12.775 1.755 12.945 8.450 ;
        RECT 17.355 1.755 17.525 8.450 ;
        RECT 21.935 1.755 22.105 8.450 ;
        RECT 26.515 1.755 26.685 8.450 ;
        RECT 31.095 1.755 31.265 8.450 ;
        RECT 35.675 1.755 35.845 8.450 ;
        RECT 40.255 1.755 40.425 8.450 ;
        RECT 44.835 1.755 45.005 8.450 ;
        RECT 49.415 1.755 49.585 8.450 ;
        RECT 53.995 1.755 54.165 8.450 ;
        RECT 58.575 1.755 58.745 8.450 ;
        RECT 63.155 1.755 63.325 8.450 ;
        RECT 67.735 1.755 67.905 8.450 ;
        RECT 72.315 1.755 72.485 8.450 ;
        RECT 76.895 1.755 77.065 8.450 ;
        RECT 81.475 1.755 81.645 8.450 ;
        RECT 86.055 1.755 86.225 8.450 ;
        RECT 90.635 1.755 90.805 8.450 ;
        RECT 95.215 1.755 95.385 8.450 ;
        RECT 99.795 1.755 99.965 8.450 ;
        RECT 104.375 1.755 104.545 8.450 ;
        RECT 108.955 1.755 109.125 8.450 ;
        RECT 113.535 1.755 113.705 8.450 ;
        RECT 118.115 1.755 118.285 8.450 ;
        RECT 122.695 1.755 122.865 8.450 ;
        RECT 127.275 1.755 127.445 8.450 ;
        RECT 131.855 1.755 132.025 8.450 ;
        RECT 136.435 1.755 136.605 8.450 ;
      LAYER mcon ;
        RECT 3.615 1.835 3.785 8.165 ;
        RECT 8.195 1.835 8.365 8.165 ;
        RECT 12.775 1.835 12.945 8.165 ;
        RECT 17.355 1.835 17.525 8.165 ;
        RECT 21.935 1.835 22.105 8.165 ;
        RECT 26.515 1.835 26.685 8.165 ;
        RECT 31.095 1.835 31.265 8.165 ;
        RECT 35.675 1.835 35.845 8.165 ;
        RECT 40.255 1.835 40.425 8.165 ;
        RECT 44.835 1.835 45.005 8.165 ;
        RECT 49.415 1.835 49.585 8.165 ;
        RECT 53.995 1.835 54.165 8.165 ;
        RECT 58.575 1.835 58.745 8.165 ;
        RECT 63.155 1.835 63.325 8.165 ;
        RECT 67.735 1.835 67.905 8.165 ;
        RECT 72.315 1.835 72.485 8.165 ;
        RECT 76.895 1.835 77.065 8.165 ;
        RECT 81.475 1.835 81.645 8.165 ;
        RECT 86.055 1.835 86.225 8.165 ;
        RECT 90.635 1.835 90.805 8.165 ;
        RECT 95.215 1.835 95.385 8.165 ;
        RECT 99.795 1.835 99.965 8.165 ;
        RECT 104.375 1.835 104.545 8.165 ;
        RECT 108.955 1.835 109.125 8.165 ;
        RECT 113.535 1.835 113.705 8.165 ;
        RECT 118.115 1.835 118.285 8.165 ;
        RECT 122.695 1.835 122.865 8.165 ;
        RECT 127.275 1.835 127.445 8.165 ;
        RECT 131.855 1.835 132.025 8.165 ;
        RECT 136.435 1.835 136.605 8.165 ;
      LAYER met1 ;
        RECT 3.585 1.775 3.815 8.225 ;
        RECT 8.165 1.775 8.395 8.225 ;
        RECT 12.745 1.775 12.975 8.225 ;
        RECT 17.325 1.775 17.555 8.225 ;
        RECT 21.905 1.775 22.135 8.225 ;
        RECT 26.485 1.775 26.715 8.225 ;
        RECT 31.065 1.775 31.295 8.225 ;
        RECT 35.645 1.775 35.875 8.225 ;
        RECT 40.225 1.775 40.455 8.225 ;
        RECT 44.805 1.775 45.035 8.225 ;
        RECT 49.385 1.775 49.615 8.225 ;
        RECT 53.965 1.775 54.195 8.225 ;
        RECT 58.545 1.775 58.775 8.225 ;
        RECT 63.125 1.775 63.355 8.225 ;
        RECT 67.705 1.775 67.935 8.225 ;
        RECT 72.285 1.775 72.515 8.225 ;
        RECT 76.865 1.775 77.095 8.225 ;
        RECT 81.445 1.775 81.675 8.225 ;
        RECT 86.025 1.775 86.255 8.225 ;
        RECT 90.605 1.775 90.835 8.225 ;
        RECT 95.185 1.775 95.415 8.225 ;
        RECT 99.765 1.775 99.995 8.225 ;
        RECT 104.345 1.775 104.575 8.225 ;
        RECT 108.925 1.775 109.155 8.225 ;
        RECT 113.505 1.775 113.735 8.225 ;
        RECT 118.085 1.775 118.315 8.225 ;
        RECT 122.665 1.775 122.895 8.225 ;
        RECT 127.245 1.775 127.475 8.225 ;
        RECT 131.825 1.775 132.055 8.225 ;
        RECT 136.405 1.775 136.635 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.350 1.495 8.245 ;
        RECT 5.905 1.350 6.075 8.245 ;
        RECT 10.485 1.350 10.655 8.245 ;
        RECT 15.065 1.350 15.235 8.245 ;
        RECT 19.645 1.350 19.815 8.245 ;
        RECT 24.225 1.350 24.395 8.245 ;
        RECT 28.805 1.350 28.975 8.245 ;
        RECT 33.385 1.350 33.555 8.245 ;
        RECT 37.965 1.350 38.135 8.245 ;
        RECT 42.545 1.350 42.715 8.245 ;
        RECT 47.125 1.350 47.295 8.245 ;
        RECT 51.705 1.350 51.875 8.245 ;
        RECT 56.285 1.350 56.455 8.245 ;
        RECT 60.865 1.350 61.035 8.245 ;
        RECT 65.445 1.350 65.615 8.245 ;
        RECT 70.025 1.350 70.195 8.245 ;
        RECT 74.605 1.350 74.775 8.245 ;
        RECT 79.185 1.350 79.355 8.245 ;
        RECT 83.765 1.350 83.935 8.245 ;
        RECT 88.345 1.350 88.515 8.245 ;
        RECT 92.925 1.350 93.095 8.245 ;
        RECT 97.505 1.350 97.675 8.245 ;
        RECT 102.085 1.350 102.255 8.245 ;
        RECT 106.665 1.350 106.835 8.245 ;
        RECT 111.245 1.350 111.415 8.245 ;
        RECT 115.825 1.350 115.995 8.245 ;
        RECT 120.405 1.350 120.575 8.245 ;
        RECT 124.985 1.350 125.155 8.245 ;
        RECT 129.565 1.350 129.735 8.245 ;
        RECT 134.145 1.350 134.315 8.245 ;
        RECT 138.725 1.350 138.895 8.245 ;
        RECT 1.090 1.050 139.130 1.350 ;
      LAYER mcon ;
        RECT 1.325 1.835 1.495 8.165 ;
        RECT 5.905 1.835 6.075 8.165 ;
        RECT 10.485 1.835 10.655 8.165 ;
        RECT 15.065 1.835 15.235 8.165 ;
        RECT 19.645 1.835 19.815 8.165 ;
        RECT 24.225 1.835 24.395 8.165 ;
        RECT 28.805 1.835 28.975 8.165 ;
        RECT 33.385 1.835 33.555 8.165 ;
        RECT 37.965 1.835 38.135 8.165 ;
        RECT 42.545 1.835 42.715 8.165 ;
        RECT 47.125 1.835 47.295 8.165 ;
        RECT 51.705 1.835 51.875 8.165 ;
        RECT 56.285 1.835 56.455 8.165 ;
        RECT 60.865 1.835 61.035 8.165 ;
        RECT 65.445 1.835 65.615 8.165 ;
        RECT 70.025 1.835 70.195 8.165 ;
        RECT 74.605 1.835 74.775 8.165 ;
        RECT 79.185 1.835 79.355 8.165 ;
        RECT 83.765 1.835 83.935 8.165 ;
        RECT 88.345 1.835 88.515 8.165 ;
        RECT 92.925 1.835 93.095 8.165 ;
        RECT 97.505 1.835 97.675 8.165 ;
        RECT 102.085 1.835 102.255 8.165 ;
        RECT 106.665 1.835 106.835 8.165 ;
        RECT 111.245 1.835 111.415 8.165 ;
        RECT 115.825 1.835 115.995 8.165 ;
        RECT 120.405 1.835 120.575 8.165 ;
        RECT 124.985 1.835 125.155 8.165 ;
        RECT 129.565 1.835 129.735 8.165 ;
        RECT 134.145 1.835 134.315 8.165 ;
        RECT 138.725 1.835 138.895 8.165 ;
      LAYER met1 ;
        RECT 1.295 1.775 1.525 8.225 ;
        RECT 5.875 1.775 6.105 8.225 ;
        RECT 10.455 1.775 10.685 8.225 ;
        RECT 15.035 1.775 15.265 8.225 ;
        RECT 19.615 1.775 19.845 8.225 ;
        RECT 24.195 1.775 24.425 8.225 ;
        RECT 28.775 1.775 29.005 8.225 ;
        RECT 33.355 1.775 33.585 8.225 ;
        RECT 37.935 1.775 38.165 8.225 ;
        RECT 42.515 1.775 42.745 8.225 ;
        RECT 47.095 1.775 47.325 8.225 ;
        RECT 51.675 1.775 51.905 8.225 ;
        RECT 56.255 1.775 56.485 8.225 ;
        RECT 60.835 1.775 61.065 8.225 ;
        RECT 65.415 1.775 65.645 8.225 ;
        RECT 69.995 1.775 70.225 8.225 ;
        RECT 74.575 1.775 74.805 8.225 ;
        RECT 79.155 1.775 79.385 8.225 ;
        RECT 83.735 1.775 83.965 8.225 ;
        RECT 88.315 1.775 88.545 8.225 ;
        RECT 92.895 1.775 93.125 8.225 ;
        RECT 97.475 1.775 97.705 8.225 ;
        RECT 102.055 1.775 102.285 8.225 ;
        RECT 106.635 1.775 106.865 8.225 ;
        RECT 111.215 1.775 111.445 8.225 ;
        RECT 115.795 1.775 116.025 8.225 ;
        RECT 120.375 1.775 120.605 8.225 ;
        RECT 124.955 1.775 125.185 8.225 ;
        RECT 129.535 1.775 129.765 8.225 ;
        RECT 134.115 1.775 134.345 8.225 ;
        RECT 138.695 1.775 138.925 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 8.535 139.130 9.700 ;
        RECT 0.600 1.470 139.135 8.535 ;
        RECT 1.085 1.465 139.135 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 139.130 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
        RECT 5.980 8.850 6.780 9.250 ;
        RECT 12.480 8.850 13.280 9.250 ;
        RECT 18.980 8.850 19.780 9.250 ;
        RECT 25.480 8.850 26.280 9.250 ;
        RECT 31.980 8.850 32.780 9.250 ;
        RECT 38.480 8.850 39.280 9.250 ;
        RECT 44.980 8.850 45.780 9.250 ;
        RECT 51.480 8.850 52.280 9.250 ;
        RECT 57.980 8.850 58.780 9.250 ;
        RECT 64.480 8.850 65.280 9.250 ;
        RECT 70.980 8.850 71.780 9.250 ;
        RECT 77.480 8.850 78.280 9.250 ;
        RECT 83.980 8.850 84.780 9.250 ;
        RECT 90.480 8.850 91.280 9.250 ;
        RECT 96.980 8.850 97.780 9.250 ;
        RECT 103.480 8.850 104.280 9.250 ;
        RECT 109.980 8.850 110.780 9.250 ;
        RECT 116.480 8.850 117.280 9.250 ;
        RECT 122.980 8.850 123.780 9.250 ;
        RECT 129.480 8.850 130.280 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
        RECT 21.940 9.250 22.240 9.550 ;
        RECT 23.940 9.250 24.240 9.550 ;
        RECT 25.940 9.250 26.240 9.550 ;
        RECT 27.940 9.250 28.240 9.550 ;
        RECT 29.940 9.250 30.240 9.550 ;
        RECT 31.940 9.250 32.240 9.550 ;
        RECT 33.940 9.250 34.240 9.550 ;
        RECT 35.940 9.250 36.240 9.550 ;
        RECT 37.940 9.250 38.240 9.550 ;
        RECT 39.940 9.250 40.240 9.550 ;
        RECT 41.940 9.250 42.240 9.550 ;
        RECT 43.940 9.250 44.240 9.550 ;
        RECT 45.940 9.250 46.240 9.550 ;
        RECT 47.940 9.250 48.240 9.550 ;
        RECT 49.940 9.250 50.240 9.550 ;
        RECT 51.940 9.250 52.240 9.550 ;
        RECT 53.940 9.250 54.240 9.550 ;
        RECT 55.940 9.250 56.240 9.550 ;
        RECT 57.940 9.250 58.240 9.550 ;
        RECT 59.940 9.250 60.240 9.550 ;
        RECT 61.940 9.250 62.240 9.550 ;
        RECT 63.940 9.250 64.240 9.550 ;
        RECT 65.940 9.250 66.240 9.550 ;
        RECT 67.940 9.250 68.240 9.550 ;
        RECT 69.940 9.250 70.240 9.550 ;
        RECT 71.940 9.250 72.240 9.550 ;
        RECT 73.940 9.250 74.240 9.550 ;
        RECT 75.940 9.250 76.240 9.550 ;
        RECT 77.940 9.250 78.240 9.550 ;
        RECT 79.940 9.250 80.240 9.550 ;
        RECT 81.940 9.250 82.240 9.550 ;
        RECT 83.940 9.250 84.240 9.550 ;
        RECT 85.940 9.250 86.240 9.550 ;
        RECT 87.940 9.250 88.240 9.550 ;
        RECT 89.940 9.250 90.240 9.550 ;
        RECT 91.940 9.250 92.240 9.550 ;
        RECT 93.940 9.250 94.240 9.550 ;
        RECT 95.940 9.250 96.240 9.550 ;
        RECT 97.940 9.250 98.240 9.550 ;
        RECT 99.940 9.250 100.240 9.550 ;
        RECT 101.940 9.250 102.240 9.550 ;
        RECT 103.940 9.250 104.240 9.550 ;
        RECT 105.940 9.250 106.240 9.550 ;
        RECT 107.940 9.250 108.240 9.550 ;
        RECT 109.940 9.250 110.240 9.550 ;
        RECT 111.940 9.250 112.240 9.550 ;
        RECT 113.940 9.250 114.240 9.550 ;
        RECT 115.940 9.250 116.240 9.550 ;
        RECT 117.940 9.250 118.240 9.550 ;
        RECT 119.940 9.250 120.240 9.550 ;
        RECT 121.940 9.250 122.240 9.550 ;
        RECT 123.940 9.250 124.240 9.550 ;
        RECT 125.940 9.250 126.240 9.550 ;
        RECT 127.940 9.250 128.240 9.550 ;
        RECT 129.940 9.250 130.240 9.550 ;
        RECT 131.940 9.250 132.240 9.550 ;
        RECT 133.940 9.250 134.240 9.550 ;
        RECT 135.940 9.250 136.240 9.550 ;
        RECT 137.940 9.250 138.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 139.130 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 139.130 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
        RECT 21.940 -0.150 22.240 0.150 ;
        RECT 23.940 -0.150 24.240 0.150 ;
        RECT 25.940 -0.150 26.240 0.150 ;
        RECT 27.940 -0.150 28.240 0.150 ;
        RECT 29.940 -0.150 30.240 0.150 ;
        RECT 31.940 -0.150 32.240 0.150 ;
        RECT 33.940 -0.150 34.240 0.150 ;
        RECT 35.940 -0.150 36.240 0.150 ;
        RECT 37.940 -0.150 38.240 0.150 ;
        RECT 39.940 -0.150 40.240 0.150 ;
        RECT 41.940 -0.150 42.240 0.150 ;
        RECT 43.940 -0.150 44.240 0.150 ;
        RECT 45.940 -0.150 46.240 0.150 ;
        RECT 47.940 -0.150 48.240 0.150 ;
        RECT 49.940 -0.150 50.240 0.150 ;
        RECT 51.940 -0.150 52.240 0.150 ;
        RECT 53.940 -0.150 54.240 0.150 ;
        RECT 55.940 -0.150 56.240 0.150 ;
        RECT 57.940 -0.150 58.240 0.150 ;
        RECT 59.940 -0.150 60.240 0.150 ;
        RECT 61.940 -0.150 62.240 0.150 ;
        RECT 63.940 -0.150 64.240 0.150 ;
        RECT 65.940 -0.150 66.240 0.150 ;
        RECT 67.940 -0.150 68.240 0.150 ;
        RECT 69.940 -0.150 70.240 0.150 ;
        RECT 71.940 -0.150 72.240 0.150 ;
        RECT 73.940 -0.150 74.240 0.150 ;
        RECT 75.940 -0.150 76.240 0.150 ;
        RECT 77.940 -0.150 78.240 0.150 ;
        RECT 79.940 -0.150 80.240 0.150 ;
        RECT 81.940 -0.150 82.240 0.150 ;
        RECT 83.940 -0.150 84.240 0.150 ;
        RECT 85.940 -0.150 86.240 0.150 ;
        RECT 87.940 -0.150 88.240 0.150 ;
        RECT 89.940 -0.150 90.240 0.150 ;
        RECT 91.940 -0.150 92.240 0.150 ;
        RECT 93.940 -0.150 94.240 0.150 ;
        RECT 95.940 -0.150 96.240 0.150 ;
        RECT 97.940 -0.150 98.240 0.150 ;
        RECT 99.940 -0.150 100.240 0.150 ;
        RECT 101.940 -0.150 102.240 0.150 ;
        RECT 103.940 -0.150 104.240 0.150 ;
        RECT 105.940 -0.150 106.240 0.150 ;
        RECT 107.940 -0.150 108.240 0.150 ;
        RECT 109.940 -0.150 110.240 0.150 ;
        RECT 111.940 -0.150 112.240 0.150 ;
        RECT 113.940 -0.150 114.240 0.150 ;
        RECT 115.940 -0.150 116.240 0.150 ;
        RECT 117.940 -0.150 118.240 0.150 ;
        RECT 119.940 -0.150 120.240 0.150 ;
        RECT 121.940 -0.150 122.240 0.150 ;
        RECT 123.940 -0.150 124.240 0.150 ;
        RECT 125.940 -0.150 126.240 0.150 ;
        RECT 127.940 -0.150 128.240 0.150 ;
        RECT 129.940 -0.150 130.240 0.150 ;
        RECT 131.940 -0.150 132.240 0.150 ;
        RECT 133.940 -0.150 134.240 0.150 ;
        RECT 135.940 -0.150 136.240 0.150 ;
        RECT 137.940 -0.150 138.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 139.130 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60

#--------EOF---------

MACRO sky130_asc_res_xhigh_po_2p85_2
  CLASS CORE ;
  FOREIGN sky130_asc_res_xhigh_po_2p85_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.470 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 0.760 5.395 2.810 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 0.760 0.595 2.810 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.710 9.100 15.770 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.140 -0.300 14.340 8.250 ;
      LAYER met1 ;
        RECT 0.710 -0.300 15.770 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.710 9.250 15.770 9.550 ;
        RECT 0.705 5.375 2.865 8.225 ;
        RECT 0.705 0.575 2.865 3.425 ;
        RECT 6.700 0.150 9.780 4.850 ;
        RECT 13.615 0.575 15.775 8.225 ;
        RECT 0.710 -0.150 15.770 0.150 ;
      LAYER mcon ;
        RECT 1.560 9.250 1.860 9.550 ;
        RECT 2.560 9.250 2.860 9.550 ;
        RECT 3.560 9.250 3.860 9.550 ;
        RECT 4.560 9.250 4.860 9.550 ;
        RECT 5.560 9.250 5.860 9.550 ;
        RECT 6.560 9.250 6.860 9.550 ;
        RECT 7.560 9.250 7.860 9.550 ;
        RECT 8.560 9.250 8.860 9.550 ;
        RECT 9.560 9.250 9.860 9.550 ;
        RECT 10.560 9.250 10.860 9.550 ;
        RECT 11.560 9.250 11.860 9.550 ;
        RECT 12.560 9.250 12.860 9.550 ;
        RECT 13.560 9.250 13.860 9.550 ;
        RECT 14.560 9.250 14.860 9.550 ;
        RECT 0.795 5.455 2.780 8.145 ;
        RECT 13.700 5.455 15.685 8.145 ;
        RECT 0.795 0.655 2.780 3.345 ;
        RECT 13.700 0.655 15.685 3.345 ;
        RECT 1.560 -0.150 1.860 0.150 ;
        RECT 2.560 -0.150 2.860 0.150 ;
        RECT 3.560 -0.150 3.860 0.150 ;
        RECT 4.560 -0.150 4.860 0.150 ;
        RECT 5.560 -0.150 5.860 0.150 ;
        RECT 6.560 -0.150 6.860 0.150 ;
        RECT 7.560 -0.150 7.860 0.150 ;
        RECT 8.560 -0.150 8.860 0.150 ;
        RECT 9.560 -0.150 9.860 0.150 ;
        RECT 10.560 -0.150 10.860 0.150 ;
        RECT 11.560 -0.150 11.860 0.150 ;
        RECT 12.560 -0.150 12.860 0.150 ;
        RECT 13.560 -0.150 13.860 0.150 ;
        RECT 14.560 -0.150 14.860 0.150 ;
      LAYER met1 ;
        RECT 13.670 5.395 15.720 8.205 ;
        RECT 13.615 0.575 15.775 5.395 ;
  END
END sky130_asc_res_xhigh_po_2p85_2

#--------EOF---------

MACRO sky130_asc_pnp_05v5_W3p40L3p40_1
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.900 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.559999 ;
    PORT
      LAYER met1 ;
        RECT 2.425 3.175 5.475 6.225 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 6.408000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 6.745 6.355 7.105 ;
        RECT 1.545 2.655 1.905 6.745 ;
        RECT 5.995 2.655 6.355 6.745 ;
        RECT 1.545 2.295 6.355 2.655 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.988700 ;
    PORT
      LAYER pwell ;
        RECT 0.600 7.285 7.300 8.050 ;
        RECT 0.600 2.115 1.365 7.285 ;
        RECT 6.535 2.115 7.300 7.285 ;
        RECT 0.600 1.350 7.300 2.115 ;
      LAYER li1 ;
        RECT 0.730 7.425 7.170 7.920 ;
        RECT 0.730 1.975 1.225 7.425 ;
        RECT 6.675 1.975 7.170 7.425 ;
        RECT 0.730 1.480 7.170 1.975 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.600 9.100 7.300 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.600 -0.300 7.300 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.600 9.250 7.300 9.550 ;
        RECT 2.215 2.965 5.685 6.435 ;
        RECT 0.600 -0.150 7.300 0.150 ;
      LAYER mcon ;
        RECT 1.450 9.250 1.750 9.550 ;
        RECT 2.450 9.250 2.750 9.550 ;
        RECT 3.450 9.250 3.750 9.550 ;
        RECT 4.450 9.250 4.750 9.550 ;
        RECT 5.450 9.250 5.750 9.550 ;
        RECT 6.450 9.250 6.750 9.550 ;
        RECT 2.580 5.830 2.750 6.000 ;
        RECT 3.080 5.830 3.250 6.000 ;
        RECT 3.580 5.830 3.750 6.000 ;
        RECT 4.080 5.830 4.250 6.000 ;
        RECT 4.580 5.830 4.750 6.000 ;
        RECT 5.080 5.830 5.250 6.000 ;
        RECT 2.580 5.330 2.750 5.500 ;
        RECT 3.080 5.330 3.250 5.500 ;
        RECT 3.580 5.330 3.750 5.500 ;
        RECT 4.080 5.330 4.250 5.500 ;
        RECT 4.580 5.330 4.750 5.500 ;
        RECT 5.080 5.330 5.250 5.500 ;
        RECT 2.580 4.830 2.750 5.000 ;
        RECT 3.080 4.830 3.250 5.000 ;
        RECT 3.580 4.830 3.750 5.000 ;
        RECT 4.080 4.830 4.250 5.000 ;
        RECT 4.580 4.830 4.750 5.000 ;
        RECT 5.080 4.830 5.250 5.000 ;
        RECT 2.580 4.330 2.750 4.500 ;
        RECT 3.080 4.330 3.250 4.500 ;
        RECT 3.580 4.330 3.750 4.500 ;
        RECT 4.080 4.330 4.250 4.500 ;
        RECT 4.580 4.330 4.750 4.500 ;
        RECT 5.080 4.330 5.250 4.500 ;
        RECT 2.580 3.830 2.750 4.000 ;
        RECT 3.080 3.830 3.250 4.000 ;
        RECT 3.580 3.830 3.750 4.000 ;
        RECT 4.080 3.830 4.250 4.000 ;
        RECT 4.580 3.830 4.750 4.000 ;
        RECT 5.080 3.830 5.250 4.000 ;
        RECT 2.580 3.330 2.750 3.500 ;
        RECT 3.080 3.330 3.250 3.500 ;
        RECT 3.580 3.330 3.750 3.500 ;
        RECT 4.080 3.330 4.250 3.500 ;
        RECT 4.580 3.330 4.750 3.500 ;
        RECT 5.080 3.330 5.250 3.500 ;
        RECT 1.450 -0.150 1.750 0.150 ;
        RECT 2.450 -0.150 2.750 0.150 ;
        RECT 3.450 -0.150 3.750 0.150 ;
        RECT 4.450 -0.150 4.750 0.150 ;
        RECT 5.450 -0.150 5.750 0.150 ;
        RECT 6.450 -0.150 6.750 0.150 ;
  END
END sky130_asc_pnp_05v5_W3p40L3p40_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_12
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.815 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 154.800003 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 29.210 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.223000 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 29.210 8.650 ;
        RECT 3.615 1.755 3.785 8.450 ;
        RECT 8.195 1.755 8.365 8.450 ;
        RECT 12.775 1.755 12.945 8.450 ;
        RECT 17.355 1.755 17.525 8.450 ;
        RECT 21.935 1.755 22.105 8.450 ;
        RECT 26.515 1.755 26.685 8.450 ;
      LAYER mcon ;
        RECT 3.615 1.835 3.785 8.165 ;
        RECT 8.195 1.835 8.365 8.165 ;
        RECT 12.775 1.835 12.945 8.165 ;
        RECT 17.355 1.835 17.525 8.165 ;
        RECT 21.935 1.835 22.105 8.165 ;
        RECT 26.515 1.835 26.685 8.165 ;
      LAYER met1 ;
        RECT 3.585 1.775 3.815 8.225 ;
        RECT 8.165 1.775 8.395 8.225 ;
        RECT 12.745 1.775 12.975 8.225 ;
        RECT 17.325 1.775 17.555 8.225 ;
        RECT 21.905 1.775 22.135 8.225 ;
        RECT 26.485 1.775 26.715 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.093500 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.350 1.495 8.245 ;
        RECT 5.905 1.350 6.075 8.245 ;
        RECT 10.485 1.350 10.655 8.245 ;
        RECT 15.065 1.350 15.235 8.245 ;
        RECT 19.645 1.350 19.815 8.245 ;
        RECT 24.225 1.350 24.395 8.245 ;
        RECT 28.805 1.350 28.975 8.245 ;
        RECT 1.090 1.050 29.210 1.350 ;
      LAYER mcon ;
        RECT 1.325 1.835 1.495 8.165 ;
        RECT 5.905 1.835 6.075 8.165 ;
        RECT 10.485 1.835 10.655 8.165 ;
        RECT 15.065 1.835 15.235 8.165 ;
        RECT 19.645 1.835 19.815 8.165 ;
        RECT 24.225 1.835 24.395 8.165 ;
        RECT 28.805 1.835 28.975 8.165 ;
      LAYER met1 ;
        RECT 1.295 1.775 1.525 8.225 ;
        RECT 5.875 1.775 6.105 8.225 ;
        RECT 10.455 1.775 10.685 8.225 ;
        RECT 15.035 1.775 15.265 8.225 ;
        RECT 19.615 1.775 19.845 8.225 ;
        RECT 24.195 1.775 24.425 8.225 ;
        RECT 28.775 1.775 29.005 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 8.535 29.210 9.700 ;
        RECT 0.600 1.470 29.215 8.535 ;
        RECT 1.085 1.465 29.215 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 29.210 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
        RECT 5.980 8.850 6.780 9.250 ;
        RECT 12.480 8.850 13.280 9.250 ;
        RECT 18.980 8.850 19.780 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
        RECT 21.940 9.250 22.240 9.550 ;
        RECT 23.940 9.250 24.240 9.550 ;
        RECT 25.940 9.250 26.240 9.550 ;
        RECT 27.940 9.250 28.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 29.210 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 29.210 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
        RECT 21.940 -0.150 22.240 0.150 ;
        RECT 23.940 -0.150 24.240 0.150 ;
        RECT 25.940 -0.150 26.240 0.150 ;
        RECT 27.940 -0.150 28.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 29.210 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_12

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.590 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 72.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.520 21.990 1.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 1.090 8.450 21.990 8.750 ;
        RECT 3.435 7.020 3.605 8.450 ;
        RECT 8.015 7.020 8.185 8.450 ;
        RECT 12.595 7.020 12.765 8.450 ;
        RECT 17.175 7.020 17.345 8.450 ;
        RECT 21.755 7.020 21.925 8.450 ;
        RECT 3.435 6.930 3.610 7.020 ;
        RECT 8.015 6.930 8.190 7.020 ;
        RECT 12.595 6.930 12.770 7.020 ;
        RECT 17.175 6.930 17.350 7.020 ;
        RECT 21.755 6.930 21.930 7.020 ;
        RECT 3.440 2.980 3.610 6.930 ;
        RECT 8.020 2.980 8.190 6.930 ;
        RECT 12.600 2.980 12.770 6.930 ;
        RECT 17.180 2.980 17.350 6.930 ;
        RECT 21.760 2.980 21.930 6.930 ;
      LAYER mcon ;
        RECT 3.440 3.060 3.610 6.940 ;
        RECT 8.020 3.060 8.190 6.940 ;
        RECT 12.600 3.060 12.770 6.940 ;
        RECT 17.180 3.060 17.350 6.940 ;
        RECT 21.760 3.060 21.930 6.940 ;
      LAYER met1 ;
        RECT 3.410 3.000 3.640 7.000 ;
        RECT 7.990 3.000 8.220 7.000 ;
        RECT 12.570 3.000 12.800 7.000 ;
        RECT 17.150 3.000 17.380 7.000 ;
        RECT 21.730 3.000 21.960 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 1.150 3.270 1.320 7.020 ;
        RECT 5.730 3.270 5.900 7.020 ;
        RECT 10.310 3.270 10.480 7.020 ;
        RECT 14.890 3.270 15.060 7.020 ;
        RECT 19.470 3.270 19.640 7.020 ;
        RECT 1.145 2.980 1.320 3.270 ;
        RECT 5.725 2.980 5.900 3.270 ;
        RECT 10.305 2.980 10.480 3.270 ;
        RECT 14.885 2.980 15.060 3.270 ;
        RECT 19.465 2.980 19.640 3.270 ;
        RECT 1.145 2.650 1.315 2.980 ;
        RECT 5.725 2.650 5.895 2.980 ;
        RECT 10.305 2.650 10.475 2.980 ;
        RECT 14.885 2.650 15.055 2.980 ;
        RECT 19.465 2.650 19.635 2.980 ;
        RECT 1.090 2.350 21.990 2.650 ;
      LAYER mcon ;
        RECT 1.150 3.060 1.320 6.940 ;
        RECT 5.730 3.060 5.900 6.940 ;
        RECT 10.310 3.060 10.480 6.940 ;
        RECT 14.890 3.060 15.060 6.940 ;
        RECT 19.470 3.060 19.640 6.940 ;
      LAYER met1 ;
        RECT 1.120 3.000 1.350 7.000 ;
        RECT 5.700 3.000 5.930 7.000 ;
        RECT 10.280 3.000 10.510 7.000 ;
        RECT 14.860 3.000 15.090 7.000 ;
        RECT 19.440 3.000 19.670 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.600 9.250 21.990 9.550 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 21.990 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.600 0.150 21.990 7.130 ;
      LAYER li1 ;
        RECT 0.740 0.150 1.040 1.200 ;
        RECT 5.990 0.150 6.790 0.750 ;
        RECT 12.490 0.150 13.290 0.750 ;
        RECT 0.600 -0.150 21.990 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 21.990 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_9

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.975 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 15.470 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 15.470 8.650 ;
        RECT 3.615 1.755 3.785 8.450 ;
        RECT 8.195 1.755 8.365 8.450 ;
        RECT 12.775 1.755 12.945 8.450 ;
      LAYER mcon ;
        RECT 3.615 1.835 3.785 8.165 ;
        RECT 8.195 1.835 8.365 8.165 ;
        RECT 12.775 1.835 12.945 8.165 ;
      LAYER met1 ;
        RECT 3.585 1.775 3.815 8.225 ;
        RECT 8.165 1.775 8.395 8.225 ;
        RECT 12.745 1.775 12.975 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.350 1.495 8.245 ;
        RECT 5.905 1.350 6.075 8.245 ;
        RECT 10.485 1.350 10.655 8.245 ;
        RECT 15.065 1.350 15.235 8.245 ;
        RECT 1.090 1.050 15.470 1.350 ;
      LAYER mcon ;
        RECT 1.325 1.835 1.495 8.165 ;
        RECT 5.905 1.835 6.075 8.165 ;
        RECT 10.485 1.835 10.655 8.165 ;
        RECT 15.065 1.835 15.235 8.165 ;
      LAYER met1 ;
        RECT 1.295 1.775 1.525 8.225 ;
        RECT 5.875 1.775 6.105 8.225 ;
        RECT 10.455 1.775 10.685 8.225 ;
        RECT 15.035 1.775 15.265 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 8.535 15.470 9.700 ;
        RECT 0.600 1.470 15.475 8.535 ;
        RECT 1.085 1.465 15.475 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 15.470 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
        RECT 5.980 8.850 6.780 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 15.470 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 15.470 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 15.470 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_6

#--------EOF---------

MACRO sky130_asc_pnp_05v5_W3p40L3p40_7
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_7 ;
  ORIGIN 0.000 0.000 ;
  SIZE 48.100 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 80.919998 ;
    PORT
      LAYER met1 ;
        RECT 2.420 3.170 45.680 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 187.102295 ;
    ANTENNADIFFAREA 44.855999 ;
    PORT
      LAYER met1 ;
        RECT 1.550 6.750 46.550 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 93.967300 ;
    PORT
      LAYER pwell ;
        RECT 0.600 7.285 47.500 8.050 ;
        RECT 0.600 2.115 1.365 7.285 ;
        RECT 6.535 2.115 8.065 7.285 ;
        RECT 13.235 2.115 14.765 7.285 ;
        RECT 19.935 2.115 21.465 7.285 ;
        RECT 26.635 2.115 28.165 7.285 ;
        RECT 33.335 2.115 34.865 7.285 ;
        RECT 40.035 2.115 41.565 7.285 ;
        RECT 46.735 2.115 47.500 7.285 ;
        RECT 0.600 1.350 47.500 2.115 ;
      LAYER met1 ;
        RECT 0.730 7.500 47.370 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.600 9.100 47.500 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.600 -0.300 47.500 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.600 9.250 47.500 9.550 ;
        RECT 0.730 7.425 47.370 7.920 ;
        RECT 0.730 1.975 1.225 7.425 ;
        RECT 1.545 6.745 6.355 7.105 ;
        RECT 1.545 2.655 1.905 6.745 ;
        RECT 2.215 2.965 5.685 6.435 ;
        RECT 5.995 2.655 6.355 6.745 ;
        RECT 1.545 2.295 6.355 2.655 ;
        RECT 6.675 1.975 7.925 7.425 ;
        RECT 8.245 6.745 13.055 7.105 ;
        RECT 8.245 2.655 8.605 6.745 ;
        RECT 8.915 2.965 12.385 6.435 ;
        RECT 12.695 2.655 13.055 6.745 ;
        RECT 8.245 2.295 13.055 2.655 ;
        RECT 13.375 1.975 14.625 7.425 ;
        RECT 14.945 6.745 19.755 7.105 ;
        RECT 14.945 2.655 15.305 6.745 ;
        RECT 15.615 2.965 19.085 6.435 ;
        RECT 19.395 2.655 19.755 6.745 ;
        RECT 14.945 2.295 19.755 2.655 ;
        RECT 20.075 1.975 21.325 7.425 ;
        RECT 21.645 6.745 26.455 7.105 ;
        RECT 21.645 2.655 22.005 6.745 ;
        RECT 22.315 2.965 25.785 6.435 ;
        RECT 26.095 2.655 26.455 6.745 ;
        RECT 21.645 2.295 26.455 2.655 ;
        RECT 26.775 1.975 28.025 7.425 ;
        RECT 28.345 6.745 33.155 7.105 ;
        RECT 28.345 2.655 28.705 6.745 ;
        RECT 29.015 2.965 32.485 6.435 ;
        RECT 32.795 2.655 33.155 6.745 ;
        RECT 28.345 2.295 33.155 2.655 ;
        RECT 33.475 1.975 34.725 7.425 ;
        RECT 35.045 6.745 39.855 7.105 ;
        RECT 35.045 2.655 35.405 6.745 ;
        RECT 35.715 2.965 39.185 6.435 ;
        RECT 39.495 2.655 39.855 6.745 ;
        RECT 35.045 2.295 39.855 2.655 ;
        RECT 40.175 1.975 41.425 7.425 ;
        RECT 41.745 6.745 46.555 7.105 ;
        RECT 41.745 2.655 42.105 6.745 ;
        RECT 42.415 2.965 45.885 6.435 ;
        RECT 46.195 2.655 46.555 6.745 ;
        RECT 41.745 2.295 46.555 2.655 ;
        RECT 46.875 1.975 47.370 7.425 ;
        RECT 0.730 1.480 47.370 1.975 ;
        RECT 0.600 -0.150 47.500 0.150 ;
      LAYER mcon ;
        RECT 1.450 9.250 1.750 9.550 ;
        RECT 2.450 9.250 2.750 9.550 ;
        RECT 3.450 9.250 3.750 9.550 ;
        RECT 4.450 9.250 4.750 9.550 ;
        RECT 5.450 9.250 5.750 9.550 ;
        RECT 6.450 9.250 6.750 9.550 ;
        RECT 7.450 9.250 7.750 9.550 ;
        RECT 8.450 9.250 8.750 9.550 ;
        RECT 9.450 9.250 9.750 9.550 ;
        RECT 10.450 9.250 10.750 9.550 ;
        RECT 11.450 9.250 11.750 9.550 ;
        RECT 12.450 9.250 12.750 9.550 ;
        RECT 13.450 9.250 13.750 9.550 ;
        RECT 14.450 9.250 14.750 9.550 ;
        RECT 15.450 9.250 15.750 9.550 ;
        RECT 16.450 9.250 16.750 9.550 ;
        RECT 17.450 9.250 17.750 9.550 ;
        RECT 18.450 9.250 18.750 9.550 ;
        RECT 19.450 9.250 19.750 9.550 ;
        RECT 20.450 9.250 20.750 9.550 ;
        RECT 21.450 9.250 21.750 9.550 ;
        RECT 22.450 9.250 22.750 9.550 ;
        RECT 23.450 9.250 23.750 9.550 ;
        RECT 24.450 9.250 24.750 9.550 ;
        RECT 25.450 9.250 25.750 9.550 ;
        RECT 26.450 9.250 26.750 9.550 ;
        RECT 27.450 9.250 27.750 9.550 ;
        RECT 28.450 9.250 28.750 9.550 ;
        RECT 29.450 9.250 29.750 9.550 ;
        RECT 30.450 9.250 30.750 9.550 ;
        RECT 31.450 9.250 31.750 9.550 ;
        RECT 32.450 9.250 32.750 9.550 ;
        RECT 33.450 9.250 33.750 9.550 ;
        RECT 34.450 9.250 34.750 9.550 ;
        RECT 35.450 9.250 35.750 9.550 ;
        RECT 36.450 9.250 36.750 9.550 ;
        RECT 37.450 9.250 37.750 9.550 ;
        RECT 38.450 9.250 38.750 9.550 ;
        RECT 39.450 9.250 39.750 9.550 ;
        RECT 40.450 9.250 40.750 9.550 ;
        RECT 41.450 9.250 41.750 9.550 ;
        RECT 42.450 9.250 42.750 9.550 ;
        RECT 43.450 9.250 43.750 9.550 ;
        RECT 44.450 9.250 44.750 9.550 ;
        RECT 45.450 9.250 45.750 9.550 ;
        RECT 46.450 9.250 46.750 9.550 ;
        RECT 0.830 7.650 1.000 7.820 ;
        RECT 1.280 7.650 1.450 7.820 ;
        RECT 1.730 7.650 1.900 7.820 ;
        RECT 2.180 7.650 2.350 7.820 ;
        RECT 2.630 7.650 2.800 7.820 ;
        RECT 3.080 7.650 3.250 7.820 ;
        RECT 3.530 7.650 3.700 7.820 ;
        RECT 3.980 7.650 4.150 7.820 ;
        RECT 4.430 7.650 4.600 7.820 ;
        RECT 4.880 7.650 5.050 7.820 ;
        RECT 5.330 7.650 5.500 7.820 ;
        RECT 5.780 7.650 5.950 7.820 ;
        RECT 6.230 7.650 6.400 7.820 ;
        RECT 6.680 7.650 6.850 7.820 ;
        RECT 7.530 7.650 7.700 7.820 ;
        RECT 7.980 7.650 8.150 7.820 ;
        RECT 8.430 7.650 8.600 7.820 ;
        RECT 8.880 7.650 9.050 7.820 ;
        RECT 9.330 7.650 9.500 7.820 ;
        RECT 9.780 7.650 9.950 7.820 ;
        RECT 10.230 7.650 10.400 7.820 ;
        RECT 10.680 7.650 10.850 7.820 ;
        RECT 11.130 7.650 11.300 7.820 ;
        RECT 11.580 7.650 11.750 7.820 ;
        RECT 12.030 7.650 12.200 7.820 ;
        RECT 12.480 7.650 12.650 7.820 ;
        RECT 12.930 7.650 13.100 7.820 ;
        RECT 13.380 7.650 13.550 7.820 ;
        RECT 14.230 7.650 14.400 7.820 ;
        RECT 14.680 7.650 14.850 7.820 ;
        RECT 15.130 7.650 15.300 7.820 ;
        RECT 15.580 7.650 15.750 7.820 ;
        RECT 16.030 7.650 16.200 7.820 ;
        RECT 16.480 7.650 16.650 7.820 ;
        RECT 16.930 7.650 17.100 7.820 ;
        RECT 17.380 7.650 17.550 7.820 ;
        RECT 17.830 7.650 18.000 7.820 ;
        RECT 18.280 7.650 18.450 7.820 ;
        RECT 18.730 7.650 18.900 7.820 ;
        RECT 19.180 7.650 19.350 7.820 ;
        RECT 19.630 7.650 19.800 7.820 ;
        RECT 20.080 7.650 20.250 7.820 ;
        RECT 20.930 7.650 21.100 7.820 ;
        RECT 21.380 7.650 21.550 7.820 ;
        RECT 21.830 7.650 22.000 7.820 ;
        RECT 22.280 7.650 22.450 7.820 ;
        RECT 22.730 7.650 22.900 7.820 ;
        RECT 23.180 7.650 23.350 7.820 ;
        RECT 23.630 7.650 23.800 7.820 ;
        RECT 24.080 7.650 24.250 7.820 ;
        RECT 24.530 7.650 24.700 7.820 ;
        RECT 24.980 7.650 25.150 7.820 ;
        RECT 25.430 7.650 25.600 7.820 ;
        RECT 25.880 7.650 26.050 7.820 ;
        RECT 26.330 7.650 26.500 7.820 ;
        RECT 26.780 7.650 26.950 7.820 ;
        RECT 27.630 7.650 27.800 7.820 ;
        RECT 28.080 7.650 28.250 7.820 ;
        RECT 28.530 7.650 28.700 7.820 ;
        RECT 28.980 7.650 29.150 7.820 ;
        RECT 29.430 7.650 29.600 7.820 ;
        RECT 29.880 7.650 30.050 7.820 ;
        RECT 30.330 7.650 30.500 7.820 ;
        RECT 30.780 7.650 30.950 7.820 ;
        RECT 31.230 7.650 31.400 7.820 ;
        RECT 31.680 7.650 31.850 7.820 ;
        RECT 32.130 7.650 32.300 7.820 ;
        RECT 32.580 7.650 32.750 7.820 ;
        RECT 33.030 7.650 33.200 7.820 ;
        RECT 33.480 7.650 33.650 7.820 ;
        RECT 34.330 7.650 34.500 7.820 ;
        RECT 34.780 7.650 34.950 7.820 ;
        RECT 35.230 7.650 35.400 7.820 ;
        RECT 35.680 7.650 35.850 7.820 ;
        RECT 36.130 7.650 36.300 7.820 ;
        RECT 36.580 7.650 36.750 7.820 ;
        RECT 37.030 7.650 37.200 7.820 ;
        RECT 37.480 7.650 37.650 7.820 ;
        RECT 37.930 7.650 38.100 7.820 ;
        RECT 38.380 7.650 38.550 7.820 ;
        RECT 38.830 7.650 39.000 7.820 ;
        RECT 39.280 7.650 39.450 7.820 ;
        RECT 39.730 7.650 39.900 7.820 ;
        RECT 40.180 7.650 40.350 7.820 ;
        RECT 41.030 7.650 41.200 7.820 ;
        RECT 41.480 7.650 41.650 7.820 ;
        RECT 41.930 7.650 42.100 7.820 ;
        RECT 42.380 7.650 42.550 7.820 ;
        RECT 42.830 7.650 43.000 7.820 ;
        RECT 43.280 7.650 43.450 7.820 ;
        RECT 43.730 7.650 43.900 7.820 ;
        RECT 44.180 7.650 44.350 7.820 ;
        RECT 44.630 7.650 44.800 7.820 ;
        RECT 45.080 7.650 45.250 7.820 ;
        RECT 45.530 7.650 45.700 7.820 ;
        RECT 45.980 7.650 46.150 7.820 ;
        RECT 46.430 7.650 46.600 7.820 ;
        RECT 46.880 7.650 47.050 7.820 ;
        RECT 1.650 6.850 1.820 7.020 ;
        RECT 2.100 6.850 2.270 7.020 ;
        RECT 2.550 6.850 2.720 7.020 ;
        RECT 3.000 6.850 3.170 7.020 ;
        RECT 3.450 6.850 3.620 7.020 ;
        RECT 3.900 6.850 4.070 7.020 ;
        RECT 4.350 6.850 4.520 7.020 ;
        RECT 4.800 6.850 4.970 7.020 ;
        RECT 5.250 6.850 5.420 7.020 ;
        RECT 5.700 6.850 5.870 7.020 ;
        RECT 6.150 6.850 6.320 7.020 ;
        RECT 2.580 5.830 2.750 6.000 ;
        RECT 3.080 5.830 3.250 6.000 ;
        RECT 3.580 5.830 3.750 6.000 ;
        RECT 4.080 5.830 4.250 6.000 ;
        RECT 4.580 5.830 4.750 6.000 ;
        RECT 5.080 5.830 5.250 6.000 ;
        RECT 2.580 5.330 2.750 5.500 ;
        RECT 3.080 5.330 3.250 5.500 ;
        RECT 3.580 5.330 3.750 5.500 ;
        RECT 4.080 5.330 4.250 5.500 ;
        RECT 4.580 5.330 4.750 5.500 ;
        RECT 5.080 5.330 5.250 5.500 ;
        RECT 2.580 4.830 2.750 5.000 ;
        RECT 3.080 4.830 3.250 5.000 ;
        RECT 3.580 4.830 3.750 5.000 ;
        RECT 4.080 4.830 4.250 5.000 ;
        RECT 4.580 4.830 4.750 5.000 ;
        RECT 5.080 4.830 5.250 5.000 ;
        RECT 2.580 4.330 2.750 4.500 ;
        RECT 3.080 4.330 3.250 4.500 ;
        RECT 3.580 4.330 3.750 4.500 ;
        RECT 4.080 4.330 4.250 4.500 ;
        RECT 4.580 4.330 4.750 4.500 ;
        RECT 5.080 4.330 5.250 4.500 ;
        RECT 2.580 3.830 2.750 4.000 ;
        RECT 3.080 3.830 3.250 4.000 ;
        RECT 3.580 3.830 3.750 4.000 ;
        RECT 4.080 3.830 4.250 4.000 ;
        RECT 4.580 3.830 4.750 4.000 ;
        RECT 5.080 3.830 5.250 4.000 ;
        RECT 2.580 3.330 2.750 3.500 ;
        RECT 3.080 3.330 3.250 3.500 ;
        RECT 3.580 3.330 3.750 3.500 ;
        RECT 4.080 3.330 4.250 3.500 ;
        RECT 4.580 3.330 4.750 3.500 ;
        RECT 5.080 3.330 5.250 3.500 ;
        RECT 8.350 6.850 8.520 7.020 ;
        RECT 8.800 6.850 8.970 7.020 ;
        RECT 9.250 6.850 9.420 7.020 ;
        RECT 9.700 6.850 9.870 7.020 ;
        RECT 10.150 6.850 10.320 7.020 ;
        RECT 10.600 6.850 10.770 7.020 ;
        RECT 11.050 6.850 11.220 7.020 ;
        RECT 11.500 6.850 11.670 7.020 ;
        RECT 11.950 6.850 12.120 7.020 ;
        RECT 12.400 6.850 12.570 7.020 ;
        RECT 12.850 6.850 13.020 7.020 ;
        RECT 9.280 5.830 9.450 6.000 ;
        RECT 9.780 5.830 9.950 6.000 ;
        RECT 10.280 5.830 10.450 6.000 ;
        RECT 10.780 5.830 10.950 6.000 ;
        RECT 11.280 5.830 11.450 6.000 ;
        RECT 11.780 5.830 11.950 6.000 ;
        RECT 9.280 5.330 9.450 5.500 ;
        RECT 9.780 5.330 9.950 5.500 ;
        RECT 10.280 5.330 10.450 5.500 ;
        RECT 10.780 5.330 10.950 5.500 ;
        RECT 11.280 5.330 11.450 5.500 ;
        RECT 11.780 5.330 11.950 5.500 ;
        RECT 9.280 4.830 9.450 5.000 ;
        RECT 9.780 4.830 9.950 5.000 ;
        RECT 10.280 4.830 10.450 5.000 ;
        RECT 10.780 4.830 10.950 5.000 ;
        RECT 11.280 4.830 11.450 5.000 ;
        RECT 11.780 4.830 11.950 5.000 ;
        RECT 9.280 4.330 9.450 4.500 ;
        RECT 9.780 4.330 9.950 4.500 ;
        RECT 10.280 4.330 10.450 4.500 ;
        RECT 10.780 4.330 10.950 4.500 ;
        RECT 11.280 4.330 11.450 4.500 ;
        RECT 11.780 4.330 11.950 4.500 ;
        RECT 9.280 3.830 9.450 4.000 ;
        RECT 9.780 3.830 9.950 4.000 ;
        RECT 10.280 3.830 10.450 4.000 ;
        RECT 10.780 3.830 10.950 4.000 ;
        RECT 11.280 3.830 11.450 4.000 ;
        RECT 11.780 3.830 11.950 4.000 ;
        RECT 9.280 3.330 9.450 3.500 ;
        RECT 9.780 3.330 9.950 3.500 ;
        RECT 10.280 3.330 10.450 3.500 ;
        RECT 10.780 3.330 10.950 3.500 ;
        RECT 11.280 3.330 11.450 3.500 ;
        RECT 11.780 3.330 11.950 3.500 ;
        RECT 15.050 6.850 15.220 7.020 ;
        RECT 15.500 6.850 15.670 7.020 ;
        RECT 15.950 6.850 16.120 7.020 ;
        RECT 16.400 6.850 16.570 7.020 ;
        RECT 16.850 6.850 17.020 7.020 ;
        RECT 17.300 6.850 17.470 7.020 ;
        RECT 17.750 6.850 17.920 7.020 ;
        RECT 18.200 6.850 18.370 7.020 ;
        RECT 18.650 6.850 18.820 7.020 ;
        RECT 19.100 6.850 19.270 7.020 ;
        RECT 19.550 6.850 19.720 7.020 ;
        RECT 15.980 5.830 16.150 6.000 ;
        RECT 16.480 5.830 16.650 6.000 ;
        RECT 16.980 5.830 17.150 6.000 ;
        RECT 17.480 5.830 17.650 6.000 ;
        RECT 17.980 5.830 18.150 6.000 ;
        RECT 18.480 5.830 18.650 6.000 ;
        RECT 15.980 5.330 16.150 5.500 ;
        RECT 16.480 5.330 16.650 5.500 ;
        RECT 16.980 5.330 17.150 5.500 ;
        RECT 17.480 5.330 17.650 5.500 ;
        RECT 17.980 5.330 18.150 5.500 ;
        RECT 18.480 5.330 18.650 5.500 ;
        RECT 15.980 4.830 16.150 5.000 ;
        RECT 16.480 4.830 16.650 5.000 ;
        RECT 16.980 4.830 17.150 5.000 ;
        RECT 17.480 4.830 17.650 5.000 ;
        RECT 17.980 4.830 18.150 5.000 ;
        RECT 18.480 4.830 18.650 5.000 ;
        RECT 15.980 4.330 16.150 4.500 ;
        RECT 16.480 4.330 16.650 4.500 ;
        RECT 16.980 4.330 17.150 4.500 ;
        RECT 17.480 4.330 17.650 4.500 ;
        RECT 17.980 4.330 18.150 4.500 ;
        RECT 18.480 4.330 18.650 4.500 ;
        RECT 15.980 3.830 16.150 4.000 ;
        RECT 16.480 3.830 16.650 4.000 ;
        RECT 16.980 3.830 17.150 4.000 ;
        RECT 17.480 3.830 17.650 4.000 ;
        RECT 17.980 3.830 18.150 4.000 ;
        RECT 18.480 3.830 18.650 4.000 ;
        RECT 15.980 3.330 16.150 3.500 ;
        RECT 16.480 3.330 16.650 3.500 ;
        RECT 16.980 3.330 17.150 3.500 ;
        RECT 17.480 3.330 17.650 3.500 ;
        RECT 17.980 3.330 18.150 3.500 ;
        RECT 18.480 3.330 18.650 3.500 ;
        RECT 21.750 6.850 21.920 7.020 ;
        RECT 22.200 6.850 22.370 7.020 ;
        RECT 22.650 6.850 22.820 7.020 ;
        RECT 23.100 6.850 23.270 7.020 ;
        RECT 23.550 6.850 23.720 7.020 ;
        RECT 24.000 6.850 24.170 7.020 ;
        RECT 24.450 6.850 24.620 7.020 ;
        RECT 24.900 6.850 25.070 7.020 ;
        RECT 25.350 6.850 25.520 7.020 ;
        RECT 25.800 6.850 25.970 7.020 ;
        RECT 26.250 6.850 26.420 7.020 ;
        RECT 22.680 5.830 22.850 6.000 ;
        RECT 23.180 5.830 23.350 6.000 ;
        RECT 23.680 5.830 23.850 6.000 ;
        RECT 24.180 5.830 24.350 6.000 ;
        RECT 24.680 5.830 24.850 6.000 ;
        RECT 25.180 5.830 25.350 6.000 ;
        RECT 22.680 5.330 22.850 5.500 ;
        RECT 23.180 5.330 23.350 5.500 ;
        RECT 23.680 5.330 23.850 5.500 ;
        RECT 24.180 5.330 24.350 5.500 ;
        RECT 24.680 5.330 24.850 5.500 ;
        RECT 25.180 5.330 25.350 5.500 ;
        RECT 22.680 4.830 22.850 5.000 ;
        RECT 23.180 4.830 23.350 5.000 ;
        RECT 23.680 4.830 23.850 5.000 ;
        RECT 24.180 4.830 24.350 5.000 ;
        RECT 24.680 4.830 24.850 5.000 ;
        RECT 25.180 4.830 25.350 5.000 ;
        RECT 22.680 4.330 22.850 4.500 ;
        RECT 23.180 4.330 23.350 4.500 ;
        RECT 23.680 4.330 23.850 4.500 ;
        RECT 24.180 4.330 24.350 4.500 ;
        RECT 24.680 4.330 24.850 4.500 ;
        RECT 25.180 4.330 25.350 4.500 ;
        RECT 22.680 3.830 22.850 4.000 ;
        RECT 23.180 3.830 23.350 4.000 ;
        RECT 23.680 3.830 23.850 4.000 ;
        RECT 24.180 3.830 24.350 4.000 ;
        RECT 24.680 3.830 24.850 4.000 ;
        RECT 25.180 3.830 25.350 4.000 ;
        RECT 22.680 3.330 22.850 3.500 ;
        RECT 23.180 3.330 23.350 3.500 ;
        RECT 23.680 3.330 23.850 3.500 ;
        RECT 24.180 3.330 24.350 3.500 ;
        RECT 24.680 3.330 24.850 3.500 ;
        RECT 25.180 3.330 25.350 3.500 ;
        RECT 28.450 6.850 28.620 7.020 ;
        RECT 28.900 6.850 29.070 7.020 ;
        RECT 29.350 6.850 29.520 7.020 ;
        RECT 29.800 6.850 29.970 7.020 ;
        RECT 30.250 6.850 30.420 7.020 ;
        RECT 30.700 6.850 30.870 7.020 ;
        RECT 31.150 6.850 31.320 7.020 ;
        RECT 31.600 6.850 31.770 7.020 ;
        RECT 32.050 6.850 32.220 7.020 ;
        RECT 32.500 6.850 32.670 7.020 ;
        RECT 32.950 6.850 33.120 7.020 ;
        RECT 29.380 5.830 29.550 6.000 ;
        RECT 29.880 5.830 30.050 6.000 ;
        RECT 30.380 5.830 30.550 6.000 ;
        RECT 30.880 5.830 31.050 6.000 ;
        RECT 31.380 5.830 31.550 6.000 ;
        RECT 31.880 5.830 32.050 6.000 ;
        RECT 29.380 5.330 29.550 5.500 ;
        RECT 29.880 5.330 30.050 5.500 ;
        RECT 30.380 5.330 30.550 5.500 ;
        RECT 30.880 5.330 31.050 5.500 ;
        RECT 31.380 5.330 31.550 5.500 ;
        RECT 31.880 5.330 32.050 5.500 ;
        RECT 29.380 4.830 29.550 5.000 ;
        RECT 29.880 4.830 30.050 5.000 ;
        RECT 30.380 4.830 30.550 5.000 ;
        RECT 30.880 4.830 31.050 5.000 ;
        RECT 31.380 4.830 31.550 5.000 ;
        RECT 31.880 4.830 32.050 5.000 ;
        RECT 29.380 4.330 29.550 4.500 ;
        RECT 29.880 4.330 30.050 4.500 ;
        RECT 30.380 4.330 30.550 4.500 ;
        RECT 30.880 4.330 31.050 4.500 ;
        RECT 31.380 4.330 31.550 4.500 ;
        RECT 31.880 4.330 32.050 4.500 ;
        RECT 29.380 3.830 29.550 4.000 ;
        RECT 29.880 3.830 30.050 4.000 ;
        RECT 30.380 3.830 30.550 4.000 ;
        RECT 30.880 3.830 31.050 4.000 ;
        RECT 31.380 3.830 31.550 4.000 ;
        RECT 31.880 3.830 32.050 4.000 ;
        RECT 29.380 3.330 29.550 3.500 ;
        RECT 29.880 3.330 30.050 3.500 ;
        RECT 30.380 3.330 30.550 3.500 ;
        RECT 30.880 3.330 31.050 3.500 ;
        RECT 31.380 3.330 31.550 3.500 ;
        RECT 31.880 3.330 32.050 3.500 ;
        RECT 35.150 6.850 35.320 7.020 ;
        RECT 35.600 6.850 35.770 7.020 ;
        RECT 36.050 6.850 36.220 7.020 ;
        RECT 36.500 6.850 36.670 7.020 ;
        RECT 36.950 6.850 37.120 7.020 ;
        RECT 37.400 6.850 37.570 7.020 ;
        RECT 37.850 6.850 38.020 7.020 ;
        RECT 38.300 6.850 38.470 7.020 ;
        RECT 38.750 6.850 38.920 7.020 ;
        RECT 39.200 6.850 39.370 7.020 ;
        RECT 39.650 6.850 39.820 7.020 ;
        RECT 36.080 5.830 36.250 6.000 ;
        RECT 36.580 5.830 36.750 6.000 ;
        RECT 37.080 5.830 37.250 6.000 ;
        RECT 37.580 5.830 37.750 6.000 ;
        RECT 38.080 5.830 38.250 6.000 ;
        RECT 38.580 5.830 38.750 6.000 ;
        RECT 36.080 5.330 36.250 5.500 ;
        RECT 36.580 5.330 36.750 5.500 ;
        RECT 37.080 5.330 37.250 5.500 ;
        RECT 37.580 5.330 37.750 5.500 ;
        RECT 38.080 5.330 38.250 5.500 ;
        RECT 38.580 5.330 38.750 5.500 ;
        RECT 36.080 4.830 36.250 5.000 ;
        RECT 36.580 4.830 36.750 5.000 ;
        RECT 37.080 4.830 37.250 5.000 ;
        RECT 37.580 4.830 37.750 5.000 ;
        RECT 38.080 4.830 38.250 5.000 ;
        RECT 38.580 4.830 38.750 5.000 ;
        RECT 36.080 4.330 36.250 4.500 ;
        RECT 36.580 4.330 36.750 4.500 ;
        RECT 37.080 4.330 37.250 4.500 ;
        RECT 37.580 4.330 37.750 4.500 ;
        RECT 38.080 4.330 38.250 4.500 ;
        RECT 38.580 4.330 38.750 4.500 ;
        RECT 36.080 3.830 36.250 4.000 ;
        RECT 36.580 3.830 36.750 4.000 ;
        RECT 37.080 3.830 37.250 4.000 ;
        RECT 37.580 3.830 37.750 4.000 ;
        RECT 38.080 3.830 38.250 4.000 ;
        RECT 38.580 3.830 38.750 4.000 ;
        RECT 36.080 3.330 36.250 3.500 ;
        RECT 36.580 3.330 36.750 3.500 ;
        RECT 37.080 3.330 37.250 3.500 ;
        RECT 37.580 3.330 37.750 3.500 ;
        RECT 38.080 3.330 38.250 3.500 ;
        RECT 38.580 3.330 38.750 3.500 ;
        RECT 41.850 6.850 42.020 7.020 ;
        RECT 42.300 6.850 42.470 7.020 ;
        RECT 42.750 6.850 42.920 7.020 ;
        RECT 43.200 6.850 43.370 7.020 ;
        RECT 43.650 6.850 43.820 7.020 ;
        RECT 44.100 6.850 44.270 7.020 ;
        RECT 44.550 6.850 44.720 7.020 ;
        RECT 45.000 6.850 45.170 7.020 ;
        RECT 45.450 6.850 45.620 7.020 ;
        RECT 45.900 6.850 46.070 7.020 ;
        RECT 46.350 6.850 46.520 7.020 ;
        RECT 42.780 5.830 42.950 6.000 ;
        RECT 43.280 5.830 43.450 6.000 ;
        RECT 43.780 5.830 43.950 6.000 ;
        RECT 44.280 5.830 44.450 6.000 ;
        RECT 44.780 5.830 44.950 6.000 ;
        RECT 45.280 5.830 45.450 6.000 ;
        RECT 42.780 5.330 42.950 5.500 ;
        RECT 43.280 5.330 43.450 5.500 ;
        RECT 43.780 5.330 43.950 5.500 ;
        RECT 44.280 5.330 44.450 5.500 ;
        RECT 44.780 5.330 44.950 5.500 ;
        RECT 45.280 5.330 45.450 5.500 ;
        RECT 42.780 4.830 42.950 5.000 ;
        RECT 43.280 4.830 43.450 5.000 ;
        RECT 43.780 4.830 43.950 5.000 ;
        RECT 44.280 4.830 44.450 5.000 ;
        RECT 44.780 4.830 44.950 5.000 ;
        RECT 45.280 4.830 45.450 5.000 ;
        RECT 42.780 4.330 42.950 4.500 ;
        RECT 43.280 4.330 43.450 4.500 ;
        RECT 43.780 4.330 43.950 4.500 ;
        RECT 44.280 4.330 44.450 4.500 ;
        RECT 44.780 4.330 44.950 4.500 ;
        RECT 45.280 4.330 45.450 4.500 ;
        RECT 42.780 3.830 42.950 4.000 ;
        RECT 43.280 3.830 43.450 4.000 ;
        RECT 43.780 3.830 43.950 4.000 ;
        RECT 44.280 3.830 44.450 4.000 ;
        RECT 44.780 3.830 44.950 4.000 ;
        RECT 45.280 3.830 45.450 4.000 ;
        RECT 42.780 3.330 42.950 3.500 ;
        RECT 43.280 3.330 43.450 3.500 ;
        RECT 43.780 3.330 43.950 3.500 ;
        RECT 44.280 3.330 44.450 3.500 ;
        RECT 44.780 3.330 44.950 3.500 ;
        RECT 45.280 3.330 45.450 3.500 ;
        RECT 1.450 -0.150 1.750 0.150 ;
        RECT 2.450 -0.150 2.750 0.150 ;
        RECT 3.450 -0.150 3.750 0.150 ;
        RECT 4.450 -0.150 4.750 0.150 ;
        RECT 5.450 -0.150 5.750 0.150 ;
        RECT 6.450 -0.150 6.750 0.150 ;
        RECT 7.450 -0.150 7.750 0.150 ;
        RECT 8.450 -0.150 8.750 0.150 ;
        RECT 9.450 -0.150 9.750 0.150 ;
        RECT 10.450 -0.150 10.750 0.150 ;
        RECT 11.450 -0.150 11.750 0.150 ;
        RECT 12.450 -0.150 12.750 0.150 ;
        RECT 13.450 -0.150 13.750 0.150 ;
        RECT 14.450 -0.150 14.750 0.150 ;
        RECT 15.450 -0.150 15.750 0.150 ;
        RECT 16.450 -0.150 16.750 0.150 ;
        RECT 17.450 -0.150 17.750 0.150 ;
        RECT 18.450 -0.150 18.750 0.150 ;
        RECT 19.450 -0.150 19.750 0.150 ;
        RECT 20.450 -0.150 20.750 0.150 ;
        RECT 21.450 -0.150 21.750 0.150 ;
        RECT 22.450 -0.150 22.750 0.150 ;
        RECT 23.450 -0.150 23.750 0.150 ;
        RECT 24.450 -0.150 24.750 0.150 ;
        RECT 25.450 -0.150 25.750 0.150 ;
        RECT 26.450 -0.150 26.750 0.150 ;
        RECT 27.450 -0.150 27.750 0.150 ;
        RECT 28.450 -0.150 28.750 0.150 ;
        RECT 29.450 -0.150 29.750 0.150 ;
        RECT 30.450 -0.150 30.750 0.150 ;
        RECT 31.450 -0.150 31.750 0.150 ;
        RECT 32.450 -0.150 32.750 0.150 ;
        RECT 33.450 -0.150 33.750 0.150 ;
        RECT 34.450 -0.150 34.750 0.150 ;
        RECT 35.450 -0.150 35.750 0.150 ;
        RECT 36.450 -0.150 36.750 0.150 ;
        RECT 37.450 -0.150 37.750 0.150 ;
        RECT 38.450 -0.150 38.750 0.150 ;
        RECT 39.450 -0.150 39.750 0.150 ;
        RECT 40.450 -0.150 40.750 0.150 ;
        RECT 41.450 -0.150 41.750 0.150 ;
        RECT 42.450 -0.150 42.750 0.150 ;
        RECT 43.450 -0.150 43.750 0.150 ;
        RECT 44.450 -0.150 44.750 0.150 ;
        RECT 45.450 -0.150 45.750 0.150 ;
        RECT 46.450 -0.150 46.750 0.150 ;
  END
END sky130_asc_pnp_05v5_W3p40L3p40_7

#--------EOF---------

MACRO sky130_asc_cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_asc_cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 37.055 BY 9.400 ;
  SITE unitasc ;
  PIN Cin
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 0.600 7.850 1.600 8.250 ;
    END
  END Cin
  PIN Cout
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 0.710 0.700 1.510 1.200 ;
    END
  END Cout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.610 9.250 36.450 9.550 ;
      LAYER mcon ;
        RECT 1.460 9.250 1.760 9.550 ;
        RECT 3.460 9.250 3.760 9.550 ;
        RECT 5.460 9.250 5.760 9.550 ;
        RECT 7.460 9.250 7.760 9.550 ;
        RECT 9.460 9.250 9.760 9.550 ;
        RECT 11.460 9.250 11.760 9.550 ;
        RECT 13.460 9.250 13.760 9.550 ;
        RECT 15.460 9.250 15.760 9.550 ;
        RECT 17.460 9.250 17.760 9.550 ;
        RECT 19.460 9.250 19.760 9.550 ;
        RECT 21.460 9.250 21.760 9.550 ;
        RECT 23.460 9.250 23.760 9.550 ;
        RECT 25.460 9.250 25.760 9.550 ;
        RECT 27.460 9.250 27.760 9.550 ;
        RECT 29.460 9.250 29.760 9.550 ;
        RECT 31.460 9.250 31.760 9.550 ;
        RECT 33.460 9.250 33.760 9.550 ;
        RECT 35.460 9.250 35.760 9.550 ;
      LAYER met1 ;
        RECT 0.610 9.100 36.450 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.610 -0.150 36.450 0.150 ;
      LAYER mcon ;
        RECT 1.460 -0.150 1.760 0.150 ;
        RECT 3.460 -0.150 3.760 0.150 ;
        RECT 5.460 -0.150 5.760 0.150 ;
        RECT 7.460 -0.150 7.760 0.150 ;
        RECT 9.460 -0.150 9.760 0.150 ;
        RECT 11.460 -0.150 11.760 0.150 ;
        RECT 13.460 -0.150 13.760 0.150 ;
        RECT 15.460 -0.150 15.760 0.150 ;
        RECT 17.460 -0.150 17.760 0.150 ;
        RECT 19.460 -0.150 19.760 0.150 ;
        RECT 21.460 -0.150 21.760 0.150 ;
        RECT 23.460 -0.150 23.760 0.150 ;
        RECT 25.460 -0.150 25.760 0.150 ;
        RECT 27.460 -0.150 27.760 0.150 ;
        RECT 29.460 -0.150 29.760 0.150 ;
        RECT 31.460 -0.150 31.760 0.150 ;
        RECT 33.460 -0.150 33.760 0.150 ;
        RECT 35.460 -0.150 35.760 0.150 ;
      LAYER met1 ;
        RECT 0.610 -0.300 36.450 0.300 ;
    END
  END VGND
  OBS
      LAYER met3 ;
        RECT 0.600 1.750 37 8.250 ;
      LAYER met4 ;
        RECT 0.4 0.500 36.830 8.870 ;
      LAYER met5 ;
        RECT 0.4 0.500 36.830 8.870 ;
  END
END sky130_asc_cap_mim_m3_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.850 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 22.350 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 22.350 8.650 ;
        RECT 3.615 8.245 3.785 8.450 ;
        RECT 8.195 8.245 8.365 8.450 ;
        RECT 12.775 8.245 12.945 8.450 ;
        RECT 17.355 8.245 17.525 8.450 ;
        RECT 21.935 8.245 22.105 8.450 ;
        RECT 3.615 8.130 3.790 8.245 ;
        RECT 8.195 8.130 8.370 8.245 ;
        RECT 12.775 8.130 12.950 8.245 ;
        RECT 17.355 8.130 17.530 8.245 ;
        RECT 21.935 8.130 22.110 8.245 ;
        RECT 3.620 1.755 3.790 8.130 ;
        RECT 8.200 1.755 8.370 8.130 ;
        RECT 12.780 1.755 12.950 8.130 ;
        RECT 17.360 1.755 17.530 8.130 ;
        RECT 21.940 1.755 22.110 8.130 ;
      LAYER mcon ;
        RECT 3.620 1.835 3.790 8.165 ;
        RECT 8.200 1.835 8.370 8.165 ;
        RECT 12.780 1.835 12.950 8.165 ;
        RECT 17.360 1.835 17.530 8.165 ;
        RECT 21.940 1.835 22.110 8.165 ;
      LAYER met1 ;
        RECT 3.590 1.775 3.820 8.225 ;
        RECT 8.170 1.775 8.400 8.225 ;
        RECT 12.750 1.775 12.980 8.225 ;
        RECT 17.330 1.775 17.560 8.225 ;
        RECT 21.910 1.775 22.140 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 1.330 1.870 1.500 8.245 ;
        RECT 5.910 1.870 6.080 8.245 ;
        RECT 10.490 1.870 10.660 8.245 ;
        RECT 15.070 1.870 15.240 8.245 ;
        RECT 19.650 1.870 19.820 8.245 ;
        RECT 1.325 1.755 1.500 1.870 ;
        RECT 5.905 1.755 6.080 1.870 ;
        RECT 10.485 1.755 10.660 1.870 ;
        RECT 15.065 1.755 15.240 1.870 ;
        RECT 19.645 1.755 19.820 1.870 ;
        RECT 1.325 1.350 1.495 1.755 ;
        RECT 5.905 1.350 6.075 1.755 ;
        RECT 10.485 1.350 10.655 1.755 ;
        RECT 15.065 1.350 15.235 1.755 ;
        RECT 19.645 1.350 19.815 1.755 ;
        RECT 1.090 1.050 22.350 1.350 ;
      LAYER mcon ;
        RECT 1.330 1.835 1.500 8.165 ;
        RECT 5.910 1.835 6.080 8.165 ;
        RECT 10.490 1.835 10.660 8.165 ;
        RECT 15.070 1.835 15.240 8.165 ;
        RECT 19.650 1.835 19.820 8.165 ;
      LAYER met1 ;
        RECT 1.300 1.775 1.530 8.225 ;
        RECT 5.880 1.775 6.110 8.225 ;
        RECT 10.460 1.775 10.690 8.225 ;
        RECT 15.040 1.775 15.270 8.225 ;
        RECT 19.620 1.775 19.850 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 1.470 22.350 9.700 ;
        RECT 1.090 1.465 22.350 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 22.350 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
        RECT 5.990 8.850 6.790 9.250 ;
        RECT 12.490 8.850 13.290 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 22.350 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 22.350 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 22.350 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9

#--------EOF---------

END LIBRARY