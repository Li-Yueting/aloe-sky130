magic
tech sky130A
magscale 1 2
timestamp 1652752851
<< nwell >>
rect 90 1707 3064 1940
rect 90 294 3065 1707
rect 187 293 3065 294
<< pmoslvt >>
rect 281 355 681 1645
rect 739 355 1139 1645
rect 1197 355 1597 1645
rect 1655 355 2055 1645
rect 2113 355 2513 1645
rect 2571 355 2971 1645
<< pdiff >>
rect 223 1633 281 1645
rect 223 367 235 1633
rect 269 367 281 1633
rect 223 355 281 367
rect 681 1633 739 1645
rect 681 367 693 1633
rect 727 367 739 1633
rect 681 355 739 367
rect 1139 1633 1197 1645
rect 1139 367 1151 1633
rect 1185 367 1197 1633
rect 1139 355 1197 367
rect 1597 1633 1655 1645
rect 1597 367 1609 1633
rect 1643 367 1655 1633
rect 1597 355 1655 367
rect 2055 1633 2113 1645
rect 2055 367 2067 1633
rect 2101 367 2113 1633
rect 2055 355 2113 367
rect 2513 1633 2571 1645
rect 2513 367 2525 1633
rect 2559 367 2571 1633
rect 2513 355 2571 367
rect 2971 1633 3029 1645
rect 2971 367 2983 1633
rect 3017 367 3029 1633
rect 2971 355 3029 367
<< pdiffc >>
rect 235 367 269 1633
rect 693 367 727 1633
rect 1151 367 1185 1633
rect 1609 367 1643 1633
rect 2067 367 2101 1633
rect 2525 367 2559 1633
rect 2983 367 3017 1633
<< nsubdiff >>
rect 128 1760 168 1800
rect 128 1680 168 1720
<< nsubdiffcont >>
rect 128 1720 168 1760
<< poly >>
rect 281 1645 681 1671
rect 739 1645 1139 1671
rect 1197 1645 1597 1671
rect 1655 1645 2055 1671
rect 2113 1645 2513 1671
rect 2571 1645 2971 1671
rect 281 329 681 355
rect 739 329 1139 355
rect 1197 329 1597 355
rect 1655 329 2055 355
rect 2113 329 2513 355
rect 2571 329 2971 355
rect 428 184 548 329
rect 884 184 1004 329
rect 1340 184 1460 329
rect 1796 184 1916 329
rect 2252 184 2372 329
rect 2708 184 2828 329
rect 188 164 3064 184
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3064 164
rect 188 84 3064 104
<< polycont >>
rect 358 104 418 164
rect 758 104 818 164
rect 1158 104 1218 164
rect 1558 104 1618 164
rect 1958 104 2018 164
rect 2358 104 2418 164
rect 2758 104 2818 164
<< locali >>
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3064 1910
rect 118 1760 178 1850
rect 118 1720 128 1760
rect 168 1720 178 1760
rect 248 1730 3064 1790
rect 118 1640 178 1720
rect 235 1633 269 1649
rect 235 270 269 367
rect 693 1633 727 1730
rect 693 351 727 367
rect 1151 1633 1185 1649
rect 1151 270 1185 367
rect 1609 1633 1643 1730
rect 1609 351 1643 367
rect 2067 1633 2101 1649
rect 2067 270 2101 367
rect 2525 1633 2559 1730
rect 2525 351 2559 367
rect 2983 1633 3017 1649
rect 2983 270 3017 367
rect 188 210 3064 270
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3064 164
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3064 30
<< viali >>
rect 358 1850 418 1910
rect 758 1850 818 1910
rect 1158 1850 1218 1910
rect 1558 1850 1618 1910
rect 1958 1850 2018 1910
rect 2358 1850 2418 1910
rect 2758 1850 2818 1910
rect 235 367 269 1633
rect 693 367 727 1633
rect 1151 367 1185 1633
rect 1609 367 1643 1633
rect 2067 367 2101 1633
rect 2525 367 2559 1633
rect 2983 367 3017 1633
rect 358 -30 418 30
rect 758 -30 818 30
rect 1158 -30 1218 30
rect 1558 -30 1618 30
rect 1958 -30 2018 30
rect 2358 -30 2418 30
rect 2758 -30 2818 30
<< metal1 >>
rect 90 1910 3064 1940
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3064 1910
rect 90 1820 3064 1850
rect 229 1633 275 1645
rect 229 367 235 1633
rect 269 367 275 1633
rect 229 355 275 367
rect 687 1633 733 1645
rect 687 367 693 1633
rect 727 367 733 1633
rect 687 355 733 367
rect 1145 1633 1191 1645
rect 1145 367 1151 1633
rect 1185 367 1191 1633
rect 1145 355 1191 367
rect 1603 1633 1649 1645
rect 1603 367 1609 1633
rect 1643 367 1649 1633
rect 1603 355 1649 367
rect 2061 1633 2107 1645
rect 2061 367 2067 1633
rect 2101 367 2107 1633
rect 2061 355 2107 367
rect 2519 1633 2565 1645
rect 2519 367 2525 1633
rect 2559 367 2565 1633
rect 2519 355 2565 367
rect 2977 1633 3023 1645
rect 2977 367 2983 1633
rect 3017 367 3023 1633
rect 2977 355 3023 367
rect 90 30 3064 60
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3064 30
rect 90 -60 3064 -30
<< labels >>
flabel nwell 90 1850 150 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 90 -30 248 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 3004 1730 3064 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 3004 210 3064 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 3004 104 3064 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3155 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
