VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.750 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 21.750 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 21.750 8.950 ;
        RECT 3.015 8.245 3.185 8.650 ;
        RECT 7.595 8.245 7.765 8.650 ;
        RECT 12.175 8.245 12.345 8.650 ;
        RECT 16.755 8.245 16.925 8.650 ;
        RECT 21.335 8.245 21.505 8.650 ;
        RECT 3.015 8.130 3.190 8.245 ;
        RECT 7.595 8.130 7.770 8.245 ;
        RECT 12.175 8.130 12.350 8.245 ;
        RECT 16.755 8.130 16.930 8.245 ;
        RECT 21.335 8.130 21.510 8.245 ;
        RECT 3.020 1.755 3.190 8.130 ;
        RECT 7.600 1.755 7.770 8.130 ;
        RECT 12.180 1.755 12.350 8.130 ;
        RECT 16.760 1.755 16.930 8.130 ;
        RECT 21.340 1.755 21.510 8.130 ;
      LAYER mcon ;
        RECT 3.020 1.835 3.190 8.165 ;
        RECT 7.600 1.835 7.770 8.165 ;
        RECT 12.180 1.835 12.350 8.165 ;
        RECT 16.760 1.835 16.930 8.165 ;
        RECT 21.340 1.835 21.510 8.165 ;
      LAYER met1 ;
        RECT 2.990 1.775 3.220 8.225 ;
        RECT 7.570 1.775 7.800 8.225 ;
        RECT 12.150 1.775 12.380 8.225 ;
        RECT 16.730 1.775 16.960 8.225 ;
        RECT 21.310 1.775 21.540 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.730 1.870 0.900 8.245 ;
        RECT 5.310 1.870 5.480 8.245 ;
        RECT 9.890 1.870 10.060 8.245 ;
        RECT 14.470 1.870 14.640 8.245 ;
        RECT 19.050 1.870 19.220 8.245 ;
        RECT 0.725 1.755 0.900 1.870 ;
        RECT 5.305 1.755 5.480 1.870 ;
        RECT 9.885 1.755 10.060 1.870 ;
        RECT 14.465 1.755 14.640 1.870 ;
        RECT 19.045 1.755 19.220 1.870 ;
        RECT 0.725 1.350 0.895 1.755 ;
        RECT 5.305 1.350 5.475 1.755 ;
        RECT 9.885 1.350 10.055 1.755 ;
        RECT 14.465 1.350 14.635 1.755 ;
        RECT 19.045 1.350 19.215 1.755 ;
        RECT 0.490 1.050 21.750 1.350 ;
      LAYER mcon ;
        RECT 0.730 1.835 0.900 8.165 ;
        RECT 5.310 1.835 5.480 8.165 ;
        RECT 9.890 1.835 10.060 8.165 ;
        RECT 14.470 1.835 14.640 8.165 ;
        RECT 19.050 1.835 19.220 8.165 ;
      LAYER met1 ;
        RECT 0.700 1.775 0.930 8.225 ;
        RECT 5.280 1.775 5.510 8.225 ;
        RECT 9.860 1.775 10.090 8.225 ;
        RECT 14.440 1.775 14.670 8.225 ;
        RECT 19.020 1.775 19.250 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.470 21.750 9.700 ;
        RECT 0.490 1.465 21.750 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 21.750 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
        RECT 15.340 9.250 15.640 9.550 ;
        RECT 17.340 9.250 17.640 9.550 ;
        RECT 19.340 9.250 19.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 21.750 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 21.750 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
        RECT 15.340 -0.150 15.640 0.150 ;
        RECT 17.340 -0.150 17.640 0.150 ;
        RECT 19.340 -0.150 19.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 21.750 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9
END LIBRARY

