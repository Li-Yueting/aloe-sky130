VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.630 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.510 3.590 0.810 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.650 8.650 3.590 8.950 ;
        RECT 3.175 8.245 3.345 8.650 ;
        RECT 3.175 8.130 3.350 8.245 ;
        RECT 3.180 1.755 3.350 8.130 ;
      LAYER mcon ;
        RECT 3.180 1.835 3.350 8.165 ;
      LAYER met1 ;
        RECT 3.150 1.775 3.380 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.890 1.860 1.060 8.245 ;
        RECT 0.885 1.755 1.060 1.860 ;
        RECT 0.885 1.350 1.055 1.755 ;
        RECT 0.650 1.050 3.590 1.350 ;
      LAYER mcon ;
        RECT 0.890 1.835 1.060 8.165 ;
      LAYER met1 ;
        RECT 0.860 1.775 1.090 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.650 9.250 3.590 9.550 ;
      LAYER mcon ;
        RECT 1.500 9.250 1.800 9.550 ;
      LAYER met1 ;
        RECT 0.650 9.100 3.590 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.650 -0.150 3.590 0.150 ;
      LAYER mcon ;
        RECT 1.500 -0.150 1.800 0.150 ;
      LAYER met1 ;
        RECT 0.650 -0.300 3.590 0.300 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.650 1.465 3.590 9.700 ;
  END
END sky130_asc_pfet_01v8_lvt_1
END LIBRARY

