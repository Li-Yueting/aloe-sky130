magic
tech sky130A
magscale 1 2
timestamp 1654756426
<< locali >>
rect 576794 586112 577600 586136
rect 576794 586008 576844 586112
rect 577304 586098 577600 586112
rect 577304 586029 577995 586098
rect 577304 586008 577600 586029
rect 576794 585974 577600 586008
rect 577604 584818 577734 584860
rect 577926 584612 577995 586029
rect 577586 584552 577995 584612
rect 577926 584548 577995 584552
rect 576802 496678 577416 496712
rect 576802 496608 576918 496678
rect 577268 496608 577416 496678
rect 577564 496635 578109 496700
rect 576802 496576 577416 496608
rect 577792 495464 577938 495474
rect 577792 495456 577814 495464
rect 577616 495418 577814 495456
rect 577792 495398 577814 495418
rect 577914 495398 577938 495464
rect 577792 495370 577938 495398
rect 578044 495210 578109 496635
rect 577596 495150 578109 495210
rect 578044 495148 578109 495150
rect 576830 452232 577448 452268
rect 576830 452142 576898 452232
rect 577348 452142 577448 452232
rect 577590 452176 578236 452240
rect 576830 452114 577448 452142
rect 577880 451006 578028 451022
rect 577880 451000 577892 451006
rect 577656 450958 577892 451000
rect 577880 450946 577892 450958
rect 578004 450946 578028 451006
rect 577880 450926 578028 450946
rect 578172 450752 578236 452176
rect 577638 450692 578236 450752
rect 578172 450690 578236 450692
rect 576788 407774 577420 407824
rect 576788 407706 576864 407774
rect 577316 407706 577420 407774
rect 577564 407737 578227 407802
rect 576788 407670 577420 407706
rect 577846 406566 578016 406590
rect 577846 406560 577866 406566
rect 577606 406518 577866 406560
rect 577846 406486 577866 406518
rect 577984 406486 578016 406566
rect 577846 406464 578016 406486
rect 578162 406312 578227 407737
rect 577588 406252 578227 406312
rect 578162 406250 578227 406252
<< viali >>
rect 576844 586008 577304 586112
rect 577734 584794 577824 584878
rect 576918 496608 577268 496678
rect 577814 495398 577914 495464
rect 576898 452142 577348 452232
rect 577892 450946 578004 451006
rect 576864 407706 577316 407774
rect 577866 406486 577984 406566
<< metal1 >>
rect 576832 586112 577316 586118
rect 576832 586008 576844 586112
rect 577304 586008 577316 586112
rect 576832 586002 577316 586008
rect 577722 584878 577836 584884
rect 577722 584794 577734 584878
rect 577824 584794 577836 584878
rect 577722 584788 577836 584794
rect 513802 577318 514204 577372
rect 513802 577092 513886 577318
rect 514202 577092 514204 577318
rect 513802 577066 514204 577092
rect 576906 496678 577280 496684
rect 576906 496608 576918 496678
rect 577268 496608 577280 496678
rect 576906 496602 577280 496608
rect 577802 495464 577926 495470
rect 577802 495398 577814 495464
rect 577914 495398 577926 495464
rect 577802 495392 577926 495398
rect 576886 452232 577360 452238
rect 576886 452142 576898 452232
rect 577348 452142 577360 452232
rect 576886 452136 577360 452142
rect 577880 451006 578016 451012
rect 577880 450946 577892 451006
rect 578004 450946 578016 451006
rect 577880 450940 578016 450946
rect 576852 407774 577328 407780
rect 576852 407706 576864 407774
rect 577316 407706 577328 407774
rect 576852 407700 577328 407706
rect 577854 406566 577996 406572
rect 577854 406486 577866 406566
rect 577984 406486 577996 406566
rect 577854 406480 577996 406486
<< via1 >>
rect 576844 586008 577304 586112
rect 577734 584794 577824 584878
rect 513886 577092 514202 577318
rect 576918 496608 577268 496678
rect 577814 495398 577914 495464
rect 576898 452142 577348 452232
rect 577892 450946 578004 451006
rect 576864 407706 577316 407774
rect 577866 406486 577984 406566
<< metal2 >>
rect 576844 586112 577304 586122
rect 576844 585998 577304 586008
rect 577734 584878 577824 584888
rect 577734 584784 577824 584794
rect 513744 577318 514296 577394
rect 513744 577092 513886 577318
rect 514202 577092 514296 577318
rect 513744 577026 514296 577092
rect 547144 553408 548282 553488
rect 547144 552942 547302 553408
rect 548128 552942 548282 553408
rect 547144 552838 548282 552942
rect 547392 544344 547594 544370
rect 547392 544258 547438 544344
rect 547568 544258 547594 544344
rect 547392 544226 547594 544258
rect 576918 496678 577268 496688
rect 576918 496598 577268 496608
rect 577814 495464 577914 495474
rect 577814 495388 577914 495398
rect 576898 452232 577348 452242
rect 576898 452132 577348 452142
rect 577892 451006 578004 451016
rect 577892 450936 578004 450946
rect 576864 407774 577316 407784
rect 576864 407696 577316 407706
rect 577866 406566 577984 406576
rect 577866 406476 577984 406486
<< via2 >>
rect 576844 586008 577304 586112
rect 577734 584794 577824 584878
rect 513886 577092 514202 577318
rect 547302 552942 548128 553408
rect 547438 544258 547568 544344
rect 576918 496608 577268 496678
rect 576898 452142 577348 452232
rect 576864 407706 577316 407774
<< metal3 >>
rect 510594 697122 515394 702340
rect 510186 697030 515954 697122
rect 520594 697072 525394 702340
rect 510186 692630 510580 697030
rect 515380 692630 515954 697030
rect 510186 692500 515954 692630
rect 520336 697000 525630 697072
rect 520336 692600 520594 697000
rect 525394 692600 525630 697000
rect 520336 692474 525630 692600
rect 566472 644568 582450 644574
rect 562478 644114 582450 644568
rect 562478 640214 562980 644114
rect 567032 640214 582450 644114
rect 562478 639796 582450 640214
rect 566472 639778 582450 639796
rect 562482 633660 582464 634554
rect 562482 630618 563210 633660
rect 566486 630618 582464 633660
rect 562482 629758 582464 630618
rect 562354 607454 567618 607626
rect 483478 607260 567618 607454
rect 483478 607252 566960 607260
rect 483478 607244 563736 607252
rect 483478 607116 562852 607244
rect 477114 600836 477124 607116
rect 483470 607052 562852 607116
rect 563052 607236 563736 607244
rect 563052 607052 563302 607236
rect 483470 607044 563302 607052
rect 563502 607044 563736 607236
rect 563944 607044 564178 607252
rect 564386 607044 564638 607252
rect 564846 607244 566960 607252
rect 564846 607044 565114 607244
rect 483470 607036 565114 607044
rect 565322 607234 566960 607244
rect 565322 607036 565564 607234
rect 483470 607026 565564 607036
rect 565772 607026 566024 607234
rect 566232 607026 566500 607234
rect 566708 607052 566960 607234
rect 567168 607052 567618 607260
rect 566708 607026 567618 607052
rect 483470 606710 567618 607026
rect 483470 606700 564204 606710
rect 483470 606492 562852 606700
rect 563060 606492 563310 606700
rect 563518 606684 564204 606700
rect 563518 606492 563752 606684
rect 483470 606476 563752 606492
rect 563960 606476 564204 606684
rect 483470 606460 564204 606476
rect 564462 606700 567618 606710
rect 564462 606692 566968 606700
rect 564462 606460 564646 606692
rect 483470 606442 564646 606460
rect 564904 606684 566016 606692
rect 564904 606442 565106 606684
rect 483470 606434 565106 606442
rect 565364 606434 565532 606684
rect 565790 606442 566016 606684
rect 566274 606442 566484 606692
rect 566742 606450 566968 606692
rect 567226 606450 567618 606700
rect 566742 606442 567618 606450
rect 565790 606434 567618 606442
rect 483470 606174 567618 606434
rect 483470 606166 563294 606174
rect 483470 605916 562852 606166
rect 563110 605924 563294 606166
rect 563552 606166 566158 606174
rect 563552 605924 563744 606166
rect 563110 605916 563744 605924
rect 564002 606158 564704 606166
rect 564002 605916 564212 606158
rect 483470 605908 564212 605916
rect 564470 605916 564704 606158
rect 564962 605916 565172 606166
rect 565430 605916 565656 606166
rect 565914 605924 566158 606166
rect 566416 606166 567618 606174
rect 566416 605924 566684 606166
rect 565914 605916 566684 605924
rect 566942 605916 567618 606166
rect 564470 605908 567618 605916
rect 483470 605598 567618 605908
rect 483470 605590 563770 605598
rect 483470 605574 563310 605590
rect 483470 605324 562842 605574
rect 563100 605340 563310 605574
rect 563568 605348 563770 605590
rect 564028 605348 564270 605598
rect 564528 605348 564780 605598
rect 565038 605590 565816 605598
rect 565038 605348 565306 605590
rect 563568 605340 565306 605348
rect 565564 605348 565816 605590
rect 566074 605590 566768 605598
rect 566074 605348 566292 605590
rect 565564 605340 566292 605348
rect 566550 605348 566768 605590
rect 567026 605348 567618 605598
rect 566550 605340 567618 605348
rect 563100 605324 567618 605340
rect 483470 605022 567618 605324
rect 483470 605014 565322 605022
rect 483470 604998 564278 605014
rect 483470 604990 563318 604998
rect 483470 604740 562834 604990
rect 563092 604748 563318 604990
rect 563576 604748 563786 604998
rect 564044 604764 564278 604998
rect 564536 604764 564772 605014
rect 565030 604772 565322 605014
rect 565580 605014 566308 605022
rect 565580 604772 565848 605014
rect 565030 604764 565848 604772
rect 566106 604772 566308 605014
rect 566566 605014 567618 605022
rect 566566 604772 566800 605014
rect 566106 604764 566800 604772
rect 567058 604764 567618 605014
rect 564044 604748 567618 604764
rect 563092 604740 567618 604748
rect 483470 604362 567618 604740
rect 483470 604346 566526 604362
rect 483470 604330 564946 604346
rect 483470 604080 562834 604330
rect 563092 604080 563352 604330
rect 563610 604080 563870 604330
rect 564128 604322 564946 604330
rect 564128 604080 564404 604322
rect 483470 604072 564404 604080
rect 564662 604096 564946 604322
rect 565204 604096 565506 604346
rect 565764 604096 566000 604346
rect 566258 604112 566526 604346
rect 566784 604112 567010 604362
rect 567268 604112 567618 604362
rect 566258 604096 567618 604112
rect 564662 604072 567618 604096
rect 483470 603644 567618 604072
rect 483470 603636 567026 603644
rect 483470 603628 564420 603636
rect 483470 603620 563862 603628
rect 483470 603612 563368 603620
rect 483470 603362 562818 603612
rect 563076 603370 563368 603612
rect 563626 603378 563862 603620
rect 564120 603386 564420 603628
rect 564678 603628 565498 603636
rect 564678 603386 564972 603628
rect 564120 603378 564972 603386
rect 565230 603386 565498 603628
rect 565756 603386 566016 603636
rect 566274 603386 566516 603636
rect 566774 603394 567026 603636
rect 567284 603394 567618 603644
rect 566774 603386 567618 603394
rect 565230 603378 567618 603386
rect 563626 603370 567618 603378
rect 563076 603362 567618 603370
rect 483470 603026 567618 603362
rect 483470 603002 567026 603026
rect 483470 602976 566550 603002
rect 483470 602960 565506 602976
rect 483470 602952 564980 602960
rect 483470 602936 564420 602952
rect 483470 602926 563368 602936
rect 483470 602676 562834 602926
rect 563092 602686 563368 602926
rect 563626 602686 563878 602936
rect 564136 602702 564420 602936
rect 564678 602710 564980 602952
rect 565238 602726 565506 602960
rect 565764 602968 566550 602976
rect 565764 602726 566024 602968
rect 565238 602718 566024 602726
rect 566282 602752 566550 602968
rect 566808 602776 567026 603002
rect 567284 602776 567618 603026
rect 566808 602752 567618 602776
rect 566282 602718 567618 602752
rect 565238 602710 567618 602718
rect 564678 602702 567618 602710
rect 564136 602686 567618 602702
rect 563092 602676 567618 602686
rect 483470 602250 567618 602676
rect 483470 602200 566066 602250
rect 483470 602184 564420 602200
rect 483470 602176 563336 602184
rect 483470 601926 562818 602176
rect 563076 601934 563336 602176
rect 563594 601934 563854 602184
rect 564112 601950 564420 602184
rect 564678 601950 565006 602200
rect 565264 601950 565524 602200
rect 565782 602000 566066 602200
rect 566324 602226 567618 602250
rect 566324 602000 566534 602226
rect 565782 601976 566534 602000
rect 566792 601976 566984 602226
rect 567242 601976 567618 602226
rect 565782 601950 567618 601976
rect 564112 601934 567618 601950
rect 563076 601926 567618 601934
rect 483470 601500 567618 601926
rect 483470 601474 564956 601500
rect 483470 601466 563886 601474
rect 483470 601458 563352 601466
rect 483470 601208 562802 601458
rect 563060 601216 563352 601458
rect 563610 601224 563886 601466
rect 564144 601224 564396 601474
rect 564654 601250 564956 601474
rect 565214 601490 567618 601500
rect 565214 601250 565532 601490
rect 564654 601240 565532 601250
rect 565790 601474 566584 601490
rect 565790 601240 566082 601474
rect 564654 601224 566082 601240
rect 566340 601240 566584 601474
rect 566842 601474 567618 601490
rect 566842 601240 567042 601474
rect 566340 601224 567042 601240
rect 567300 601224 567618 601474
rect 563610 601216 567618 601224
rect 563060 601208 567618 601216
rect 483470 600836 567618 601208
rect 483478 600788 567618 600836
rect 562354 600514 567618 600788
rect 576834 586112 577314 586117
rect 576834 586008 576844 586112
rect 577304 586008 577314 586112
rect 576834 586003 577314 586008
rect 577724 584880 577834 584883
rect 577700 584878 577880 584880
rect 577700 584794 577734 584878
rect 577824 584794 577880 584878
rect 577700 584032 577880 584794
rect 510000 583852 583688 584032
rect 510000 583312 513488 583852
rect 514146 583312 583688 583852
rect 510000 583242 583688 583312
rect 513744 577340 514296 577394
rect 513744 577140 513814 577340
rect 514030 577318 514296 577340
rect 513744 577092 513886 577140
rect 514202 577092 514296 577318
rect 513744 577026 514296 577092
rect 572580 576308 578098 577088
rect 546676 576248 578098 576308
rect 546676 576112 573008 576248
rect 546676 574916 546908 576112
rect 547420 574916 573008 576112
rect 546676 574676 573008 574916
rect 572580 574432 573008 574676
rect 577036 574432 578098 576248
rect 483722 574092 490892 574190
rect 481644 571878 481654 574092
rect 484004 573682 490892 574092
rect 484004 572370 490738 573682
rect 491694 572370 491704 573682
rect 572580 573404 578098 574432
rect 484004 571878 490892 572370
rect 483722 571786 490892 571878
rect 547106 553534 551394 553802
rect 547106 553408 550120 553534
rect 547106 552942 547302 553408
rect 548128 552942 550120 553408
rect 547106 552600 550120 552942
rect 551016 552600 551394 553534
rect 547106 552458 551394 552600
rect 547290 544572 555842 544688
rect 547290 544344 554616 544572
rect 547290 544258 547438 544344
rect 547568 544258 554616 544344
rect 547290 543922 554616 544258
rect 555754 543922 555842 544572
rect 547290 543892 555842 543922
rect 483722 523666 491024 523924
rect 482172 522000 482182 523666
rect 484144 523558 491024 523666
rect 484144 522330 490382 523558
rect 491590 522330 491600 523558
rect 484144 522000 491024 522330
rect 483722 521854 491024 522000
rect 547550 521130 577000 521304
rect 546930 519822 546940 521130
rect 548224 520942 577000 521130
rect 548224 519960 572904 520942
rect 576342 519960 577000 520942
rect 548224 519822 577000 519960
rect 547550 519672 577000 519822
rect 506108 517760 507248 518964
rect 506108 517644 506182 517760
rect 506172 516896 506182 517644
rect 507134 517644 507248 517760
rect 507134 516896 507144 517644
rect 562090 503840 568202 504092
rect 483620 503632 568202 503840
rect 477576 497422 477586 503632
rect 484462 503360 568202 503632
rect 484462 497780 562754 503360
rect 566906 497780 568202 503360
rect 484462 497422 568202 497780
rect 483620 497174 568202 497422
rect 562090 496452 568202 497174
rect 576908 496678 577278 496683
rect 576908 496608 576918 496678
rect 577268 496608 577278 496678
rect 576908 496603 577278 496608
rect 577764 494542 577976 495482
rect 514358 494536 583900 494542
rect 505298 494432 583900 494536
rect 505298 493868 506134 494432
rect 507170 493868 583900 494432
rect 505298 493776 583900 493868
rect 514358 493752 583900 493776
rect 576888 452232 577358 452237
rect 576888 452142 576898 452232
rect 577348 452142 577358 452232
rect 576888 452137 577358 452142
rect 577862 450196 578066 451024
rect 554200 450080 583840 450196
rect 554200 449506 554676 450080
rect 555748 449506 583840 450080
rect 554200 449406 583840 449506
rect 576854 407774 577326 407779
rect 576854 407706 576864 407774
rect 577316 407706 577326 407774
rect 576854 407701 577326 407706
rect 577838 405712 578104 406596
rect 543944 405612 583854 405712
rect 543944 405034 550022 405612
rect 551408 405034 583854 405612
rect 543944 404922 583854 405034
rect 543944 404920 559164 404922
<< via3 >>
rect 510580 692630 515380 697030
rect 520594 692600 525394 697000
rect 562980 640214 567032 644114
rect 563210 630618 566486 633660
rect 477124 600836 483470 607116
rect 562852 607052 563052 607244
rect 563302 607044 563502 607236
rect 563736 607044 563944 607252
rect 564178 607044 564386 607252
rect 564638 607044 564846 607252
rect 565114 607036 565322 607244
rect 565564 607026 565772 607234
rect 566024 607026 566232 607234
rect 566500 607026 566708 607234
rect 566960 607052 567168 607260
rect 562852 606492 563060 606700
rect 563310 606492 563518 606700
rect 563752 606476 563960 606684
rect 564204 606460 564462 606710
rect 564646 606442 564904 606692
rect 565106 606434 565364 606684
rect 565532 606434 565790 606684
rect 566016 606442 566274 606692
rect 566484 606442 566742 606692
rect 566968 606450 567226 606700
rect 562852 605916 563110 606166
rect 563294 605924 563552 606174
rect 563744 605916 564002 606166
rect 564212 605908 564470 606158
rect 564704 605916 564962 606166
rect 565172 605916 565430 606166
rect 565656 605916 565914 606166
rect 566158 605924 566416 606174
rect 566684 605916 566942 606166
rect 562842 605324 563100 605574
rect 563310 605340 563568 605590
rect 563770 605348 564028 605598
rect 564270 605348 564528 605598
rect 564780 605348 565038 605598
rect 565306 605340 565564 605590
rect 565816 605348 566074 605598
rect 566292 605340 566550 605590
rect 566768 605348 567026 605598
rect 562834 604740 563092 604990
rect 563318 604748 563576 604998
rect 563786 604748 564044 604998
rect 564278 604764 564536 605014
rect 564772 604764 565030 605014
rect 565322 604772 565580 605022
rect 565848 604764 566106 605014
rect 566308 604772 566566 605022
rect 566800 604764 567058 605014
rect 562834 604080 563092 604330
rect 563352 604080 563610 604330
rect 563870 604080 564128 604330
rect 564404 604072 564662 604322
rect 564946 604096 565204 604346
rect 565506 604096 565764 604346
rect 566000 604096 566258 604346
rect 566526 604112 566784 604362
rect 567010 604112 567268 604362
rect 562818 603362 563076 603612
rect 563368 603370 563626 603620
rect 563862 603378 564120 603628
rect 564420 603386 564678 603636
rect 564972 603378 565230 603628
rect 565498 603386 565756 603636
rect 566016 603386 566274 603636
rect 566516 603386 566774 603636
rect 567026 603394 567284 603644
rect 562834 602676 563092 602926
rect 563368 602686 563626 602936
rect 563878 602686 564136 602936
rect 564420 602702 564678 602952
rect 564980 602710 565238 602960
rect 565506 602726 565764 602976
rect 566024 602718 566282 602968
rect 566550 602752 566808 603002
rect 567026 602776 567284 603026
rect 562818 601926 563076 602176
rect 563336 601934 563594 602184
rect 563854 601934 564112 602184
rect 564420 601950 564678 602200
rect 565006 601950 565264 602200
rect 565524 601950 565782 602200
rect 566066 602000 566324 602250
rect 566534 601976 566792 602226
rect 566984 601976 567242 602226
rect 562802 601208 563060 601458
rect 563352 601216 563610 601466
rect 563886 601224 564144 601474
rect 564396 601224 564654 601474
rect 564956 601250 565214 601500
rect 565532 601240 565790 601490
rect 566082 601224 566340 601474
rect 566584 601240 566842 601490
rect 567042 601224 567300 601474
rect 576844 586008 577304 586112
rect 513488 583312 514146 583852
rect 513814 577318 514030 577340
rect 513814 577140 513886 577318
rect 513886 577140 514030 577318
rect 546908 574916 547420 576112
rect 573008 574432 577036 576248
rect 481654 571878 484004 574092
rect 490738 572370 491694 573682
rect 550120 552600 551016 553534
rect 554616 543922 555754 544572
rect 482182 522000 484144 523666
rect 490382 522330 491590 523558
rect 546940 519822 548224 521130
rect 572904 519960 576342 520942
rect 506182 516896 507134 517760
rect 477586 497422 484462 503632
rect 562754 497780 566906 503360
rect 576918 496608 577268 496678
rect 506134 493868 507170 494432
rect 576898 452142 577348 452232
rect 554676 449506 555748 450080
rect 576864 407706 577316 407774
rect 550022 405034 551408 405612
<< metal4 >>
rect 115026 697030 577478 697194
rect 115026 692630 510580 697030
rect 515380 697000 577478 697030
rect 515380 692630 520594 697000
rect 115026 692600 520594 692630
rect 525394 696948 577478 697000
rect 525394 696712 572774 696948
rect 573010 696712 573600 696948
rect 574000 696712 574400 696948
rect 574800 696712 575200 696948
rect 575600 696712 576000 696948
rect 576400 696712 576800 696948
rect 577200 696712 577478 696948
rect 525394 696590 577478 696712
rect 525394 696560 576000 696590
rect 525394 696300 573600 696560
rect 574000 696300 574400 696560
rect 574800 696300 575200 696560
rect 575600 696330 576000 696560
rect 576400 696528 577478 696590
rect 576400 696330 576802 696528
rect 575600 696300 576802 696330
rect 525394 696268 576802 696300
rect 577202 696268 577478 696528
rect 525394 696144 577478 696268
rect 525394 696136 575988 696144
rect 525394 696128 575204 696136
rect 525394 696112 574402 696128
rect 525394 695852 573616 696112
rect 574016 695868 574402 696112
rect 574802 695876 575204 696128
rect 575604 695884 575988 696136
rect 576388 696136 577478 696144
rect 576388 695884 576798 696136
rect 575604 695876 576798 695884
rect 577198 695876 577478 696136
rect 574802 695868 577478 695876
rect 574016 695852 577478 695868
rect 525394 695686 577478 695852
rect 525394 695678 574410 695686
rect 525394 695418 573616 695678
rect 574016 695426 574410 695678
rect 574810 695426 575186 695686
rect 575586 695426 575988 695686
rect 576388 695426 576790 695686
rect 577190 695426 577478 695686
rect 574016 695418 577478 695426
rect 525394 695184 577478 695418
rect 525394 695176 575980 695184
rect 525394 695168 575194 695176
rect 525394 694908 573616 695168
rect 574016 694908 574410 695168
rect 574810 694916 575194 695168
rect 575594 694924 575980 695176
rect 576380 695176 577478 695184
rect 576380 694924 576798 695176
rect 575594 694916 576798 694924
rect 577198 694916 577478 695176
rect 574810 694908 577478 694916
rect 525394 694676 577478 694908
rect 525394 694658 576004 694676
rect 525394 694650 575194 694658
rect 525394 694390 573616 694650
rect 574016 694390 574418 694650
rect 574818 694398 575194 694650
rect 575594 694416 576004 694658
rect 576404 694416 576814 694676
rect 577214 694416 577478 694676
rect 575594 694398 577478 694416
rect 574818 694390 577478 694398
rect 525394 694116 577478 694390
rect 525394 694108 576822 694116
rect 525394 694098 576004 694108
rect 525394 694090 574418 694098
rect 525394 693830 573616 694090
rect 574016 693838 574418 694090
rect 574818 693838 575212 694098
rect 575612 693848 576004 694098
rect 576404 693856 576822 694108
rect 577222 693856 577478 694116
rect 576404 693848 577478 693856
rect 575612 693838 577478 693848
rect 574016 693830 577478 693838
rect 525394 693582 577478 693830
rect 525394 693564 576832 693582
rect 525394 693556 576014 693564
rect 525394 693296 573616 693556
rect 574016 693548 576014 693556
rect 574016 693532 575228 693548
rect 574016 693296 574418 693532
rect 525394 693272 574418 693296
rect 574818 693288 575228 693532
rect 575628 693304 576014 693548
rect 576414 693322 576832 693564
rect 577232 693322 577478 693582
rect 576414 693304 577478 693322
rect 575628 693288 577478 693304
rect 574818 693272 577478 693288
rect 525394 693046 577478 693272
rect 525394 693038 576840 693046
rect 525394 693022 574418 693038
rect 525394 692762 573616 693022
rect 574016 692778 574418 693022
rect 574818 693030 576840 693038
rect 574818 692778 575204 693030
rect 574016 692770 575204 692778
rect 575604 692770 576022 693030
rect 576422 692786 576840 693030
rect 577240 692786 577478 693046
rect 576422 692770 577478 692786
rect 574016 692762 577478 692770
rect 525394 692600 577478 692762
rect 115026 692456 577478 692600
rect 562478 644114 567434 644568
rect 562478 640214 562980 644114
rect 567032 640214 567434 644114
rect 562478 639796 567434 640214
rect 562748 633660 567016 634224
rect 562748 630618 563210 633660
rect 566486 630618 567016 633660
rect 562748 630122 567016 630618
rect 476924 607176 483704 607448
rect 562138 607260 568034 607776
rect 562138 607252 566960 607260
rect 562138 607244 563736 607252
rect 476898 607116 483714 607176
rect 476898 600836 477124 607116
rect 483470 600836 483714 607116
rect 476898 574093 483714 600836
rect 562138 607052 562852 607244
rect 563052 607236 563736 607244
rect 563052 607052 563302 607236
rect 562138 607044 563302 607052
rect 563502 607044 563736 607236
rect 563944 607044 564178 607252
rect 564386 607044 564638 607252
rect 564846 607244 566960 607252
rect 564846 607044 565114 607244
rect 562138 607036 565114 607044
rect 565322 607234 566960 607244
rect 565322 607036 565564 607234
rect 562138 607026 565564 607036
rect 565772 607026 566024 607234
rect 566232 607026 566500 607234
rect 566708 607052 566960 607234
rect 567168 607052 568034 607260
rect 566708 607026 568034 607052
rect 562138 607010 564438 607026
rect 562138 606760 563076 607010
rect 563334 606760 563520 607010
rect 563778 606760 563986 607010
rect 564244 606776 564438 607010
rect 564696 607018 568034 607026
rect 564696 606776 564896 607018
rect 564244 606768 564896 606776
rect 565154 607010 568034 607018
rect 565154 606768 565382 607010
rect 564244 606760 565382 606768
rect 565640 606760 568034 607010
rect 562138 606710 568034 606760
rect 562138 606700 564204 606710
rect 562138 606492 562852 606700
rect 563060 606500 563310 606700
rect 563518 606684 564204 606700
rect 563518 606500 563752 606684
rect 563960 606500 564204 606684
rect 564462 606700 568034 606710
rect 564462 606692 566968 606700
rect 564462 606500 564646 606692
rect 564904 606684 566016 606692
rect 564904 606500 565106 606684
rect 565364 606500 565532 606684
rect 565790 606500 566016 606684
rect 566274 606500 566484 606692
rect 566742 606500 566968 606692
rect 567226 606500 568034 606700
rect 562138 606166 562876 606492
rect 562138 605916 562852 606166
rect 562138 605574 562876 605916
rect 562138 605324 562842 605574
rect 562138 604990 562876 605324
rect 562138 604740 562834 604990
rect 562138 604330 562876 604740
rect 567252 604362 568034 606500
rect 562138 604080 562834 604330
rect 562138 603612 562876 604080
rect 567268 604112 568034 604362
rect 567252 603644 568034 604112
rect 562138 603362 562818 603612
rect 567284 603394 568034 603644
rect 562138 602926 562876 603362
rect 567252 603026 568034 603394
rect 562138 602676 562834 602926
rect 567284 602776 568034 603026
rect 562138 602176 562876 602676
rect 562138 601926 562818 602176
rect 562138 601458 562876 601926
rect 562138 601208 562802 601458
rect 567252 601474 568034 602776
rect 567300 601224 568034 601474
rect 562138 601074 562876 601208
rect 567252 601074 568034 601224
rect 562138 600316 568034 601074
rect 576843 586112 577305 586113
rect 576843 586008 576844 586112
rect 577304 586008 577305 586112
rect 576843 586007 577305 586008
rect 513404 583852 514214 584158
rect 513404 583312 513488 583852
rect 514146 583312 514214 583852
rect 513404 577340 514214 583312
rect 513404 577140 513814 577340
rect 514030 577140 514214 577340
rect 513404 577060 514214 577140
rect 572700 576248 577824 576796
rect 546907 576112 547421 576113
rect 546907 574916 546908 576112
rect 547420 574916 547421 576112
rect 546907 574915 547421 574916
rect 572700 574432 573008 576248
rect 577036 574432 577824 576248
rect 476898 574092 484005 574093
rect 476898 571878 481654 574092
rect 484004 571878 484005 574092
rect 572700 573882 577824 574432
rect 490884 573683 490974 573860
rect 490737 573682 491695 573683
rect 490737 572370 490738 573682
rect 491694 572370 491695 573682
rect 490737 572369 491695 572370
rect 490884 572228 490974 572369
rect 476898 571877 484005 571878
rect 476898 523752 483714 571877
rect 549906 553534 551608 554566
rect 549906 552600 550120 553534
rect 551016 552600 551608 553534
rect 476898 523667 483722 523752
rect 476898 523666 484145 523667
rect 476898 522000 482182 523666
rect 484144 522000 484145 523666
rect 490381 523558 491591 523559
rect 490381 522330 490382 523558
rect 491590 522330 491591 523558
rect 490381 522329 491591 522330
rect 476898 521999 484145 522000
rect 476898 503633 483714 521999
rect 546939 521130 548225 521131
rect 546939 519822 546940 521130
rect 548224 519822 548225 521130
rect 546939 519821 548225 519822
rect 506058 517760 507280 517846
rect 506058 516896 506182 517760
rect 507134 516896 507280 517760
rect 476898 503632 484463 503633
rect 476898 497422 477586 503632
rect 484462 497422 484463 503632
rect 476898 497421 484463 497422
rect 476898 497206 483714 497421
rect 506058 494432 507280 516896
rect 506058 493868 506134 494432
rect 507170 493868 507280 494432
rect 506058 493546 507280 493868
rect 549906 405612 551608 552600
rect 554476 544572 555922 545818
rect 554476 543922 554616 544572
rect 555754 543922 555922 544572
rect 554476 450080 555922 543922
rect 571956 521538 577816 521960
rect 571956 520942 573676 521538
rect 576202 520942 577816 521538
rect 571956 519960 572904 520942
rect 576342 519960 577816 520942
rect 571956 519188 573676 519960
rect 576202 519188 577816 519960
rect 571956 519012 577816 519188
rect 561824 503360 568600 504424
rect 561824 497780 562754 503360
rect 566906 503062 568600 503360
rect 561824 497482 563152 497780
rect 567304 497482 568600 503062
rect 561824 496186 568600 497482
rect 576917 496678 577269 496679
rect 576917 496608 576918 496678
rect 577268 496608 577269 496678
rect 576917 496607 577269 496608
rect 576897 452232 577349 452233
rect 576897 452142 576898 452232
rect 577348 452142 577349 452232
rect 576897 452141 577349 452142
rect 554476 449506 554676 450080
rect 555748 449506 555922 450080
rect 554476 448700 555922 449506
rect 576863 407774 577317 407775
rect 576863 407706 576864 407774
rect 577316 407706 577317 407774
rect 576863 407705 577317 407706
rect 549906 405034 550022 405612
rect 551408 405034 551608 405612
rect 549906 404358 551608 405034
<< via4 >>
rect 572774 696712 573010 696948
rect 573600 696712 574000 696948
rect 574400 696712 574800 696948
rect 575200 696712 575600 696948
rect 576000 696712 576400 696948
rect 576800 696712 577200 696948
rect 573600 696300 574000 696560
rect 574400 696300 574800 696560
rect 575200 696300 575600 696560
rect 576000 696330 576400 696590
rect 576802 696268 577202 696528
rect 573616 695852 574016 696112
rect 574402 695868 574802 696128
rect 575204 695876 575604 696136
rect 575988 695884 576388 696144
rect 576798 695876 577198 696136
rect 573616 695418 574016 695678
rect 574410 695426 574810 695686
rect 575186 695426 575586 695686
rect 575988 695426 576388 695686
rect 576790 695426 577190 695686
rect 573616 694908 574016 695168
rect 574410 694908 574810 695168
rect 575194 694916 575594 695176
rect 575980 694924 576380 695184
rect 576798 694916 577198 695176
rect 573616 694390 574016 694650
rect 574418 694390 574818 694650
rect 575194 694398 575594 694658
rect 576004 694416 576404 694676
rect 576814 694416 577214 694676
rect 573616 693830 574016 694090
rect 574418 693838 574818 694098
rect 575212 693838 575612 694098
rect 576004 693848 576404 694108
rect 576822 693856 577222 694116
rect 573616 693296 574016 693556
rect 574418 693272 574818 693532
rect 575228 693288 575628 693548
rect 576014 693304 576414 693564
rect 576832 693322 577232 693582
rect 573616 692762 574016 693022
rect 574418 692778 574818 693038
rect 575204 692770 575604 693030
rect 576022 692770 576422 693030
rect 576840 692786 577240 693046
rect 562980 640214 567032 644114
rect 563210 630618 566486 633660
rect 563076 606760 563334 607010
rect 563520 606760 563778 607010
rect 563986 606760 564244 607010
rect 564438 606776 564696 607026
rect 564896 606768 565154 607018
rect 565382 606760 565640 607010
rect 562876 606492 563060 606500
rect 563060 606492 563310 606500
rect 563310 606492 563518 606500
rect 563518 606492 563752 606500
rect 562876 606476 563752 606492
rect 563752 606476 563960 606500
rect 563960 606476 564204 606500
rect 562876 606460 564204 606476
rect 564204 606460 564462 606500
rect 564462 606460 564646 606500
rect 562876 606442 564646 606460
rect 564646 606442 564904 606500
rect 564904 606442 565106 606500
rect 562876 606434 565106 606442
rect 565106 606434 565364 606500
rect 565364 606434 565532 606500
rect 565532 606434 565790 606500
rect 565790 606442 566016 606500
rect 566016 606442 566274 606500
rect 566274 606442 566484 606500
rect 566484 606442 566742 606500
rect 566742 606450 566968 606500
rect 566968 606450 567226 606500
rect 567226 606450 567252 606500
rect 566742 606442 567252 606450
rect 565790 606434 567252 606442
rect 562876 606174 567252 606434
rect 562876 606166 563294 606174
rect 562876 605916 563110 606166
rect 563110 605924 563294 606166
rect 563294 605924 563552 606174
rect 563552 606166 566158 606174
rect 563552 605924 563744 606166
rect 563110 605916 563744 605924
rect 563744 605916 564002 606166
rect 564002 606158 564704 606166
rect 564002 605916 564212 606158
rect 562876 605908 564212 605916
rect 564212 605908 564470 606158
rect 564470 605916 564704 606158
rect 564704 605916 564962 606166
rect 564962 605916 565172 606166
rect 565172 605916 565430 606166
rect 565430 605916 565656 606166
rect 565656 605916 565914 606166
rect 565914 605924 566158 606166
rect 566158 605924 566416 606174
rect 566416 606166 567252 606174
rect 566416 605924 566684 606166
rect 565914 605916 566684 605924
rect 566684 605916 566942 606166
rect 566942 605916 567252 606166
rect 564470 605908 567252 605916
rect 562876 605598 567252 605908
rect 562876 605590 563770 605598
rect 562876 605574 563310 605590
rect 562876 605324 563100 605574
rect 563100 605340 563310 605574
rect 563310 605340 563568 605590
rect 563568 605348 563770 605590
rect 563770 605348 564028 605598
rect 564028 605348 564270 605598
rect 564270 605348 564528 605598
rect 564528 605348 564780 605598
rect 564780 605348 565038 605598
rect 565038 605590 565816 605598
rect 565038 605348 565306 605590
rect 563568 605340 565306 605348
rect 565306 605340 565564 605590
rect 565564 605348 565816 605590
rect 565816 605348 566074 605598
rect 566074 605590 566768 605598
rect 566074 605348 566292 605590
rect 565564 605340 566292 605348
rect 566292 605340 566550 605590
rect 566550 605348 566768 605590
rect 566768 605348 567026 605598
rect 567026 605348 567252 605598
rect 566550 605340 567252 605348
rect 563100 605324 567252 605340
rect 562876 605022 567252 605324
rect 562876 605014 565322 605022
rect 562876 604998 564278 605014
rect 562876 604990 563318 604998
rect 562876 604740 563092 604990
rect 563092 604748 563318 604990
rect 563318 604748 563576 604998
rect 563576 604748 563786 604998
rect 563786 604748 564044 604998
rect 564044 604764 564278 604998
rect 564278 604764 564536 605014
rect 564536 604764 564772 605014
rect 564772 604764 565030 605014
rect 565030 604772 565322 605014
rect 565322 604772 565580 605022
rect 565580 605014 566308 605022
rect 565580 604772 565848 605014
rect 565030 604764 565848 604772
rect 565848 604764 566106 605014
rect 566106 604772 566308 605014
rect 566308 604772 566566 605022
rect 566566 605014 567252 605022
rect 566566 604772 566800 605014
rect 566106 604764 566800 604772
rect 566800 604764 567058 605014
rect 567058 604764 567252 605014
rect 564044 604748 567252 604764
rect 563092 604740 567252 604748
rect 562876 604362 567252 604740
rect 562876 604346 566526 604362
rect 562876 604330 564946 604346
rect 562876 604080 563092 604330
rect 563092 604080 563352 604330
rect 563352 604080 563610 604330
rect 563610 604080 563870 604330
rect 563870 604080 564128 604330
rect 564128 604322 564946 604330
rect 564128 604080 564404 604322
rect 562876 604072 564404 604080
rect 564404 604072 564662 604322
rect 564662 604096 564946 604322
rect 564946 604096 565204 604346
rect 565204 604096 565506 604346
rect 565506 604096 565764 604346
rect 565764 604096 566000 604346
rect 566000 604096 566258 604346
rect 566258 604112 566526 604346
rect 566526 604112 566784 604362
rect 566784 604112 567010 604362
rect 567010 604112 567252 604362
rect 566258 604096 567252 604112
rect 564662 604072 567252 604096
rect 562876 603644 567252 604072
rect 562876 603636 567026 603644
rect 562876 603628 564420 603636
rect 562876 603620 563862 603628
rect 562876 603612 563368 603620
rect 562876 603362 563076 603612
rect 563076 603370 563368 603612
rect 563368 603370 563626 603620
rect 563626 603378 563862 603620
rect 563862 603378 564120 603628
rect 564120 603386 564420 603628
rect 564420 603386 564678 603636
rect 564678 603628 565498 603636
rect 564678 603386 564972 603628
rect 564120 603378 564972 603386
rect 564972 603378 565230 603628
rect 565230 603386 565498 603628
rect 565498 603386 565756 603636
rect 565756 603386 566016 603636
rect 566016 603386 566274 603636
rect 566274 603386 566516 603636
rect 566516 603386 566774 603636
rect 566774 603394 567026 603636
rect 567026 603394 567252 603644
rect 566774 603386 567252 603394
rect 565230 603378 567252 603386
rect 563626 603370 567252 603378
rect 563076 603362 567252 603370
rect 562876 603026 567252 603362
rect 562876 603002 567026 603026
rect 562876 602976 566550 603002
rect 562876 602960 565506 602976
rect 562876 602952 564980 602960
rect 562876 602936 564420 602952
rect 562876 602926 563368 602936
rect 562876 602676 563092 602926
rect 563092 602686 563368 602926
rect 563368 602686 563626 602936
rect 563626 602686 563878 602936
rect 563878 602686 564136 602936
rect 564136 602702 564420 602936
rect 564420 602702 564678 602952
rect 564678 602710 564980 602952
rect 564980 602710 565238 602960
rect 565238 602726 565506 602960
rect 565506 602726 565764 602976
rect 565764 602968 566550 602976
rect 565764 602726 566024 602968
rect 565238 602718 566024 602726
rect 566024 602718 566282 602968
rect 566282 602752 566550 602968
rect 566550 602752 566808 603002
rect 566808 602776 567026 603002
rect 567026 602776 567252 603026
rect 566808 602752 567252 602776
rect 566282 602718 567252 602752
rect 565238 602710 567252 602718
rect 564678 602702 567252 602710
rect 564136 602686 567252 602702
rect 563092 602676 567252 602686
rect 562876 602250 567252 602676
rect 562876 602200 566066 602250
rect 562876 602184 564420 602200
rect 562876 602176 563336 602184
rect 562876 601926 563076 602176
rect 563076 601934 563336 602176
rect 563336 601934 563594 602184
rect 563594 601934 563854 602184
rect 563854 601934 564112 602184
rect 564112 601950 564420 602184
rect 564420 601950 564678 602200
rect 564678 601950 565006 602200
rect 565006 601950 565264 602200
rect 565264 601950 565524 602200
rect 565524 601950 565782 602200
rect 565782 602000 566066 602200
rect 566066 602000 566324 602250
rect 566324 602226 567252 602250
rect 566324 602000 566534 602226
rect 565782 601976 566534 602000
rect 566534 601976 566792 602226
rect 566792 601976 566984 602226
rect 566984 601976 567242 602226
rect 567242 601976 567252 602226
rect 565782 601950 567252 601976
rect 564112 601934 567252 601950
rect 563076 601926 567252 601934
rect 562876 601500 567252 601926
rect 562876 601474 564956 601500
rect 562876 601466 563886 601474
rect 562876 601458 563352 601466
rect 562876 601208 563060 601458
rect 563060 601216 563352 601458
rect 563352 601216 563610 601466
rect 563610 601224 563886 601466
rect 563886 601224 564144 601474
rect 564144 601224 564396 601474
rect 564396 601224 564654 601474
rect 564654 601250 564956 601474
rect 564956 601250 565214 601500
rect 565214 601490 567252 601500
rect 565214 601250 565532 601490
rect 564654 601240 565532 601250
rect 565532 601240 565790 601490
rect 565790 601474 566584 601490
rect 565790 601240 566082 601474
rect 564654 601224 566082 601240
rect 566082 601224 566340 601474
rect 566340 601240 566584 601474
rect 566584 601240 566842 601490
rect 566842 601474 567252 601490
rect 566842 601240 567042 601474
rect 566340 601224 567042 601240
rect 567042 601224 567252 601474
rect 563610 601216 567252 601224
rect 563060 601208 567252 601216
rect 562876 601074 567252 601208
rect 573166 575004 576452 576020
rect 573676 520942 576202 521538
rect 573676 519960 576202 520942
rect 573676 519188 576202 519960
rect 563152 497780 566906 503062
rect 566906 497780 567304 503062
rect 563152 497482 567304 497780
<< metal5 >>
rect 572566 696948 577476 697016
rect 572566 696712 572774 696948
rect 573010 696712 573600 696948
rect 574000 696712 574400 696948
rect 574800 696712 575200 696948
rect 575600 696712 576000 696948
rect 576400 696712 576800 696948
rect 577200 696712 577476 696948
rect 572566 696590 577476 696712
rect 572566 696560 576000 696590
rect 572566 696300 573600 696560
rect 574000 696300 574400 696560
rect 574800 696300 575200 696560
rect 575600 696330 576000 696560
rect 576400 696528 577476 696590
rect 576400 696330 576802 696528
rect 575600 696300 576802 696330
rect 572566 696268 576802 696300
rect 577202 696268 577476 696528
rect 572566 696144 577476 696268
rect 572566 696136 575988 696144
rect 572566 696128 575204 696136
rect 572566 696112 574402 696128
rect 572566 695852 573616 696112
rect 574016 695868 574402 696112
rect 574802 695876 575204 696128
rect 575604 695884 575988 696136
rect 576388 696136 577476 696144
rect 576388 695884 576798 696136
rect 575604 695876 576798 695884
rect 577198 695876 577476 696136
rect 574802 695868 577476 695876
rect 574016 695852 577476 695868
rect 572566 695686 577476 695852
rect 572566 695678 574410 695686
rect 572566 695418 573616 695678
rect 574016 695426 574410 695678
rect 574810 695426 575186 695686
rect 575586 695426 575988 695686
rect 576388 695426 576790 695686
rect 577190 695426 577476 695686
rect 574016 695418 577476 695426
rect 572566 695184 577476 695418
rect 572566 695176 575980 695184
rect 572566 695168 575194 695176
rect 572566 694908 573616 695168
rect 574016 694908 574410 695168
rect 574810 694916 575194 695168
rect 575594 694924 575980 695176
rect 576380 695176 577476 695184
rect 576380 694924 576798 695176
rect 575594 694916 576798 694924
rect 577198 694916 577476 695176
rect 574810 694908 577476 694916
rect 572566 694676 577476 694908
rect 572566 694658 576004 694676
rect 572566 694650 575194 694658
rect 572566 694390 573616 694650
rect 574016 694390 574418 694650
rect 574818 694398 575194 694650
rect 575594 694416 576004 694658
rect 576404 694416 576814 694676
rect 577214 694416 577476 694676
rect 575594 694398 577476 694416
rect 574818 694390 577476 694398
rect 572566 694116 577476 694390
rect 572566 694108 576822 694116
rect 572566 694098 576004 694108
rect 572566 694090 574418 694098
rect 572566 693830 573616 694090
rect 574016 693838 574418 694090
rect 574818 693838 575212 694098
rect 575612 693848 576004 694098
rect 576404 693856 576822 694108
rect 577222 693856 577476 694116
rect 576404 693848 577476 693856
rect 575612 693838 577476 693848
rect 574016 693830 577476 693838
rect 572566 693582 577476 693830
rect 572566 693564 576832 693582
rect 572566 693556 576014 693564
rect 572566 693296 573616 693556
rect 574016 693548 576014 693556
rect 574016 693532 575228 693548
rect 574016 693296 574418 693532
rect 572566 693272 574418 693296
rect 574818 693288 575228 693532
rect 575628 693304 576014 693548
rect 576414 693322 576832 693564
rect 577232 693322 577476 693582
rect 576414 693304 577476 693322
rect 575628 693288 577476 693304
rect 574818 693272 577476 693288
rect 572566 693046 577476 693272
rect 572566 693038 576840 693046
rect 572566 693022 574418 693038
rect 572566 692762 573616 693022
rect 574016 692778 574418 693022
rect 574818 693030 576840 693038
rect 574818 692778 575204 693030
rect 574016 692770 575204 692778
rect 575604 692770 576022 693030
rect 576422 692786 576840 693030
rect 577240 692786 577476 693046
rect 576422 692770 577476 692786
rect 574016 692762 577476 692770
rect 572566 692660 577476 692762
rect 562482 644114 567446 646728
rect 562482 640214 562980 644114
rect 567032 640214 567446 644114
rect 562482 633660 567446 640214
rect 562482 630618 563210 633660
rect 566486 630618 567446 633660
rect 562482 629784 567446 630618
rect 562456 629294 567446 629784
rect 562456 607026 567424 629294
rect 562456 607010 564438 607026
rect 562456 606760 563076 607010
rect 563334 606760 563520 607010
rect 563778 606760 563986 607010
rect 564244 606776 564438 607010
rect 564696 607018 567424 607026
rect 564696 606776 564896 607018
rect 564244 606768 564896 606776
rect 565154 607010 567424 607018
rect 565154 606768 565382 607010
rect 564244 606760 565382 606768
rect 565640 606760 567424 607010
rect 562456 606500 567424 606760
rect 562456 601074 562876 606500
rect 567252 601074 567424 606500
rect 562456 503062 567424 601074
rect 562456 497482 563152 503062
rect 567304 497482 567424 503062
rect 562456 480000 567424 497482
rect 572560 576020 577480 692660
rect 572560 575004 573166 576020
rect 576452 575004 577480 576020
rect 572560 521538 577480 575004
rect 572560 519188 573676 521538
rect 576202 519188 577480 521538
rect 572560 495782 577480 519188
rect 572562 398674 577478 495782
use bgr_top_flat  bgr_top_flat_0
timestamp 1654684494
transform 0 -1 547550 1 0 518772
box 0 0 58512 56576
use nmos_flat  nmos_flat_0
timestamp 1654747070
transform 1 0 575038 0 1 585348
box -2706 -1060 2609 940
use nmos_flat  nmos_flat_1
timestamp 1654747070
transform 1 0 575048 0 1 495946
box -2706 -1060 2609 940
use nmos_flat  nmos_flat_2
timestamp 1654747070
transform 1 0 575090 0 1 451488
box -2706 -1060 2609 940
use nmos_flat  nmos_flat_3
timestamp 1654747070
transform 1 0 575040 0 1 407048
box -2706 -1060 2609 940
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0
timestamp 1632839657
transform 1 0 0 0 1 0
box -800 -800 584800 704800
<< end >>
