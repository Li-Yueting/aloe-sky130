VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO box
  CLASS CORE ;
  FOREIGN box ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.470 BY 4.700 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.820 2.940 1.120 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.950 2.940 9.250 ;
        RECT 2.525 8.545 2.695 8.950 ;
        RECT 2.525 8.430 2.700 8.545 ;
        RECT 2.530 2.055 2.700 8.430 ;
      LAYER mcon ;
        RECT 2.530 2.135 2.700 8.465 ;
      LAYER met1 ;
        RECT 2.500 2.075 2.730 8.525 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.240 2.170 0.410 8.545 ;
        RECT 0.235 2.055 0.410 2.170 ;
        RECT 0.235 1.650 0.405 2.055 ;
        RECT 0.000 1.350 2.940 1.650 ;
      LAYER mcon ;
        RECT 0.240 2.135 0.410 8.465 ;
      LAYER met1 ;
        RECT 0.210 2.075 0.440 8.525 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.765 2.940 10.000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.550 2.940 9.850 ;
      LAYER mcon ;
        RECT 0.850 9.550 1.150 9.850 ;
      LAYER met1 ;
        RECT 0.000 9.400 2.940 10.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.150 2.940 0.450 ;
      LAYER mcon ;
        RECT 0.850 0.150 1.150 0.450 ;
      LAYER met1 ;
        RECT 0.000 0.000 2.940 0.600 ;
    END
  END VGND
END box
END LIBRARY

