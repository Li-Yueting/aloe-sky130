magic
tech sky130A
magscale 1 2
timestamp 1652142564
<< pwell >>
rect 288 -60 2728 1650
<< psubdiff >>
rect 1200 940 1816 970
rect 1200 820 1260 940
rect 1756 820 1816 940
rect 1200 790 1816 820
<< psubdiffcont >>
rect 1260 820 1756 940
<< xpolycontact >>
rect 1 1075 433 1645
rect 2583 1075 3015 1645
rect 1 115 433 685
rect 2583 115 3015 685
<< xpolyres >>
rect 433 1075 2583 1645
rect 433 115 2583 685
<< locali >>
rect 2 1850 172 1910
rect 232 1850 372 1910
rect 432 1850 572 1910
rect 632 1850 772 1910
rect 832 1850 972 1910
rect 1032 1850 1172 1910
rect 1232 1850 1372 1910
rect 1432 1850 1572 1910
rect 1632 1850 1772 1910
rect 1832 1850 1972 1910
rect 2032 1850 2172 1910
rect 2232 1850 2372 1910
rect 2432 1850 2572 1910
rect 2632 1850 2772 1910
rect 2832 1850 3014 1910
rect 1200 940 1816 970
rect 1200 820 1260 940
rect 1756 820 1816 940
rect 1200 30 1816 820
rect 2583 685 3015 1075
rect 2 -30 172 30
rect 232 -30 372 30
rect 432 -30 572 30
rect 632 -30 772 30
rect 832 -30 972 30
rect 1032 -30 1172 30
rect 1232 -30 1372 30
rect 1432 -30 1572 30
rect 1632 -30 1772 30
rect 1832 -30 1972 30
rect 2032 -30 2172 30
rect 2232 -30 2372 30
rect 2432 -30 2572 30
rect 2632 -30 2772 30
rect 2832 -30 3014 30
<< viali >>
rect 172 1850 232 1910
rect 372 1850 432 1910
rect 572 1850 632 1910
rect 772 1850 832 1910
rect 972 1850 1032 1910
rect 1172 1850 1232 1910
rect 1372 1850 1432 1910
rect 1572 1850 1632 1910
rect 1772 1850 1832 1910
rect 1972 1850 2032 1910
rect 2172 1850 2232 1910
rect 2372 1850 2432 1910
rect 2572 1850 2632 1910
rect 2772 1850 2832 1910
rect 19 1091 416 1629
rect 2600 1091 2997 1629
rect 19 131 416 669
rect 2600 131 2997 669
rect 172 -30 232 30
rect 372 -30 432 30
rect 572 -30 632 30
rect 772 -30 832 30
rect 972 -30 1032 30
rect 1172 -30 1232 30
rect 1372 -30 1432 30
rect 1572 -30 1632 30
rect 1772 -30 1832 30
rect 1972 -30 2032 30
rect 2172 -30 2232 30
rect 2372 -30 2432 30
rect 2572 -30 2632 30
rect 2772 -30 2832 30
<< metal1 >>
rect 2 1910 3014 1940
rect 2 1850 172 1910
rect 232 1850 372 1910
rect 432 1850 572 1910
rect 632 1850 772 1910
rect 832 1850 972 1910
rect 1032 1850 1172 1910
rect 1232 1850 1372 1910
rect 1432 1850 1572 1910
rect 1632 1850 1772 1910
rect 1832 1850 1972 1910
rect 2032 1850 2172 1910
rect 2232 1850 2372 1910
rect 2432 1850 2572 1910
rect 2632 1850 2772 1910
rect 2832 1850 3014 1910
rect 2 1820 3014 1850
rect 12 1629 422 1641
rect 12 1091 19 1629
rect 416 1091 422 1629
rect 12 1079 422 1091
rect 2594 1629 3004 1641
rect 2594 1091 2600 1629
rect 2997 1091 3004 1629
rect 2594 1079 3004 1091
rect 12 669 422 681
rect 12 131 19 669
rect 416 131 422 669
rect 12 119 422 131
rect 2583 669 3015 1079
rect 2583 131 2600 669
rect 2997 131 3015 669
rect 2583 115 3015 131
rect 2 30 3014 60
rect 2 -30 172 30
rect 232 -30 372 30
rect 432 -30 572 30
rect 632 -30 772 30
rect 832 -30 972 30
rect 1032 -30 1172 30
rect 1232 -30 1372 30
rect 1432 -30 1572 30
rect 1632 -30 1772 30
rect 1832 -30 1972 30
rect 2032 -30 2172 30
rect 2232 -30 2372 30
rect 2432 -30 2572 30
rect 2632 -30 2772 30
rect 2832 -30 3014 30
rect 2 -60 3014 -30
<< labels >>
flabel metal1 121 1300 241 1420 1 FreeSans 480 0 0 0 Rin
port 1 n default bidirectional
flabel metal1 121 340 241 460 1 FreeSans 480 0 0 0 Rout
port 2 n default bidirectional
flabel metal1 2 1850 62 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 2 -30 62 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 3014 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
