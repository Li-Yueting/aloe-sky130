magic
tech sky130A
magscale 1 2
timestamp 1652936965
<< nwell >>
rect 90 1707 5812 1940
rect 90 294 5813 1707
rect 187 293 5813 294
<< pmoslvt >>
rect 281 355 681 1645
rect 739 355 1139 1645
rect 1197 355 1597 1645
rect 1655 355 2055 1645
rect 2113 355 2513 1645
rect 2571 355 2971 1645
rect 3029 355 3429 1645
rect 3487 355 3887 1645
rect 3945 355 4345 1645
rect 4403 355 4803 1645
rect 4861 355 5261 1645
rect 5319 355 5719 1645
<< pdiff >>
rect 223 1633 281 1645
rect 223 367 235 1633
rect 269 367 281 1633
rect 223 355 281 367
rect 681 1633 739 1645
rect 681 367 693 1633
rect 727 367 739 1633
rect 681 355 739 367
rect 1139 1633 1197 1645
rect 1139 367 1151 1633
rect 1185 367 1197 1633
rect 1139 355 1197 367
rect 1597 1633 1655 1645
rect 1597 367 1609 1633
rect 1643 367 1655 1633
rect 1597 355 1655 367
rect 2055 1633 2113 1645
rect 2055 367 2067 1633
rect 2101 367 2113 1633
rect 2055 355 2113 367
rect 2513 1633 2571 1645
rect 2513 367 2525 1633
rect 2559 367 2571 1633
rect 2513 355 2571 367
rect 2971 1633 3029 1645
rect 2971 367 2983 1633
rect 3017 367 3029 1633
rect 2971 355 3029 367
rect 3429 1633 3487 1645
rect 3429 367 3441 1633
rect 3475 367 3487 1633
rect 3429 355 3487 367
rect 3887 1633 3945 1645
rect 3887 367 3899 1633
rect 3933 367 3945 1633
rect 3887 355 3945 367
rect 4345 1633 4403 1645
rect 4345 367 4357 1633
rect 4391 367 4403 1633
rect 4345 355 4403 367
rect 4803 1633 4861 1645
rect 4803 367 4815 1633
rect 4849 367 4861 1633
rect 4803 355 4861 367
rect 5261 1633 5319 1645
rect 5261 367 5273 1633
rect 5307 367 5319 1633
rect 5261 355 5319 367
rect 5719 1633 5777 1645
rect 5719 367 5731 1633
rect 5765 367 5777 1633
rect 5719 355 5777 367
<< pdiffc >>
rect 235 367 269 1633
rect 693 367 727 1633
rect 1151 367 1185 1633
rect 1609 367 1643 1633
rect 2067 367 2101 1633
rect 2525 367 2559 1633
rect 2983 367 3017 1633
rect 3441 367 3475 1633
rect 3899 367 3933 1633
rect 4357 367 4391 1633
rect 4815 367 4849 1633
rect 5273 367 5307 1633
rect 5731 367 5765 1633
<< nsubdiff >>
rect 1186 1808 1306 1810
rect 128 1760 168 1800
rect 1186 1772 1226 1808
rect 1270 1772 1306 1808
rect 1186 1770 1306 1772
rect 2486 1808 2606 1810
rect 2486 1772 2526 1808
rect 2570 1772 2606 1808
rect 2486 1770 2606 1772
rect 3786 1808 3906 1810
rect 3786 1772 3826 1808
rect 3870 1772 3906 1808
rect 3786 1770 3906 1772
rect 128 1680 168 1720
<< nsubdiffcont >>
rect 1226 1772 1270 1808
rect 2526 1772 2570 1808
rect 3826 1772 3870 1808
rect 128 1720 168 1760
<< poly >>
rect 281 1645 681 1671
rect 739 1645 1139 1671
rect 1197 1645 1597 1671
rect 1655 1645 2055 1671
rect 2113 1645 2513 1671
rect 2571 1645 2971 1671
rect 3029 1645 3429 1671
rect 3487 1645 3887 1671
rect 3945 1645 4345 1671
rect 4403 1645 4803 1671
rect 4861 1645 5261 1671
rect 5319 1645 5719 1671
rect 281 329 681 355
rect 739 329 1139 355
rect 1197 329 1597 355
rect 1655 329 2055 355
rect 2113 329 2513 355
rect 2571 329 2971 355
rect 3029 329 3429 355
rect 3487 329 3887 355
rect 3945 329 4345 355
rect 4403 329 4803 355
rect 4861 329 5261 355
rect 5319 329 5719 355
rect 428 184 548 329
rect 884 184 1004 329
rect 1340 184 1460 329
rect 1796 184 1916 329
rect 2252 184 2372 329
rect 2708 184 2828 329
rect 3164 184 3284 329
rect 3620 184 3740 329
rect 4076 184 4196 329
rect 4532 184 4652 329
rect 4988 184 5108 329
rect 5444 184 5564 329
rect 188 164 5812 184
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3158 164
rect 3218 104 3558 164
rect 3618 104 3958 164
rect 4018 104 4358 164
rect 4418 104 4758 164
rect 4818 104 5158 164
rect 5218 104 5558 164
rect 5618 104 5812 164
rect 188 84 5812 104
<< polycont >>
rect 358 104 418 164
rect 758 104 818 164
rect 1158 104 1218 164
rect 1558 104 1618 164
rect 1958 104 2018 164
rect 2358 104 2418 164
rect 2758 104 2818 164
rect 3158 104 3218 164
rect 3558 104 3618 164
rect 3958 104 4018 164
rect 4358 104 4418 164
rect 4758 104 4818 164
rect 5158 104 5218 164
rect 5558 104 5618 164
<< locali >>
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4358 1910
rect 4418 1850 4758 1910
rect 4818 1850 5158 1910
rect 5218 1850 5558 1910
rect 5618 1850 5812 1910
rect 118 1760 178 1850
rect 1166 1808 1326 1850
rect 1166 1772 1226 1808
rect 1270 1772 1326 1808
rect 1166 1770 1326 1772
rect 2466 1808 2626 1850
rect 2466 1772 2526 1808
rect 2570 1772 2626 1808
rect 2466 1770 2626 1772
rect 3766 1808 3926 1850
rect 3766 1772 3826 1808
rect 3870 1772 3926 1808
rect 3766 1770 3926 1772
rect 118 1720 128 1760
rect 168 1720 178 1760
rect 118 1640 178 1720
rect 248 1690 5812 1730
rect 235 1633 269 1649
rect 235 270 269 367
rect 693 1633 727 1690
rect 693 351 727 367
rect 1151 1633 1185 1649
rect 1151 270 1185 367
rect 1609 1633 1643 1690
rect 1609 351 1643 367
rect 2067 1633 2101 1649
rect 2067 270 2101 367
rect 2525 1633 2559 1690
rect 2525 351 2559 367
rect 2983 1633 3017 1649
rect 2983 270 3017 367
rect 3441 1633 3475 1690
rect 3441 351 3475 367
rect 3899 1633 3933 1649
rect 3899 270 3933 367
rect 4357 1633 4391 1690
rect 4357 351 4391 367
rect 4815 1633 4849 1649
rect 4815 270 4849 367
rect 5273 1633 5307 1690
rect 5273 351 5307 367
rect 5731 1633 5765 1649
rect 5731 270 5765 367
rect 188 210 5812 270
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3158 164
rect 3218 104 3558 164
rect 3618 104 3958 164
rect 4018 104 4358 164
rect 4418 104 4758 164
rect 4818 104 5158 164
rect 5218 104 5558 164
rect 5618 104 5812 164
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4358 30
rect 4418 -30 4758 30
rect 4818 -30 5158 30
rect 5218 -30 5558 30
rect 5618 -30 5812 30
<< viali >>
rect 358 1850 418 1910
rect 758 1850 818 1910
rect 1158 1850 1218 1910
rect 1558 1850 1618 1910
rect 1958 1850 2018 1910
rect 2358 1850 2418 1910
rect 2758 1850 2818 1910
rect 3158 1850 3218 1910
rect 3558 1850 3618 1910
rect 3958 1850 4018 1910
rect 4358 1850 4418 1910
rect 4758 1850 4818 1910
rect 5158 1850 5218 1910
rect 5558 1850 5618 1910
rect 235 367 269 1633
rect 693 367 727 1633
rect 1151 367 1185 1633
rect 1609 367 1643 1633
rect 2067 367 2101 1633
rect 2525 367 2559 1633
rect 2983 367 3017 1633
rect 3441 367 3475 1633
rect 3899 367 3933 1633
rect 4357 367 4391 1633
rect 4815 367 4849 1633
rect 5273 367 5307 1633
rect 5731 367 5765 1633
rect 358 -30 418 30
rect 758 -30 818 30
rect 1158 -30 1218 30
rect 1558 -30 1618 30
rect 1958 -30 2018 30
rect 2358 -30 2418 30
rect 2758 -30 2818 30
rect 3158 -30 3218 30
rect 3558 -30 3618 30
rect 3958 -30 4018 30
rect 4358 -30 4418 30
rect 4758 -30 4818 30
rect 5158 -30 5218 30
rect 5558 -30 5618 30
<< metal1 >>
rect 90 1910 5812 1940
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4358 1910
rect 4418 1850 4758 1910
rect 4818 1850 5158 1910
rect 5218 1850 5558 1910
rect 5618 1850 5812 1910
rect 90 1820 5812 1850
rect 229 1633 275 1645
rect 229 367 235 1633
rect 269 367 275 1633
rect 229 355 275 367
rect 687 1633 733 1645
rect 687 367 693 1633
rect 727 367 733 1633
rect 687 355 733 367
rect 1145 1633 1191 1645
rect 1145 367 1151 1633
rect 1185 367 1191 1633
rect 1145 355 1191 367
rect 1603 1633 1649 1645
rect 1603 367 1609 1633
rect 1643 367 1649 1633
rect 1603 355 1649 367
rect 2061 1633 2107 1645
rect 2061 367 2067 1633
rect 2101 367 2107 1633
rect 2061 355 2107 367
rect 2519 1633 2565 1645
rect 2519 367 2525 1633
rect 2559 367 2565 1633
rect 2519 355 2565 367
rect 2977 1633 3023 1645
rect 2977 367 2983 1633
rect 3017 367 3023 1633
rect 2977 355 3023 367
rect 3435 1633 3481 1645
rect 3435 367 3441 1633
rect 3475 367 3481 1633
rect 3435 355 3481 367
rect 3893 1633 3939 1645
rect 3893 367 3899 1633
rect 3933 367 3939 1633
rect 3893 355 3939 367
rect 4351 1633 4397 1645
rect 4351 367 4357 1633
rect 4391 367 4397 1633
rect 4351 355 4397 367
rect 4809 1633 4855 1645
rect 4809 367 4815 1633
rect 4849 367 4855 1633
rect 4809 355 4855 367
rect 5267 1633 5313 1645
rect 5267 367 5273 1633
rect 5307 367 5313 1633
rect 5267 355 5313 367
rect 5725 1633 5771 1645
rect 5725 367 5731 1633
rect 5765 367 5771 1633
rect 5725 355 5771 367
rect 90 30 5812 60
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4358 30
rect 4418 -30 4758 30
rect 4818 -30 5158 30
rect 5218 -30 5558 30
rect 5618 -30 5812 30
rect 90 -60 5812 -30
<< labels >>
flabel nwell 90 1850 150 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 90 -30 248 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 5752 1690 5812 1730 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 5752 210 5812 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 5752 104 5812 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5903 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
