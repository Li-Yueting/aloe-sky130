VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.650 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 22.200 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 22.200 8.650 ;
        RECT 3.465 8.245 3.635 8.450 ;
        RECT 8.045 8.245 8.215 8.450 ;
        RECT 12.625 8.245 12.795 8.450 ;
        RECT 17.205 8.245 17.375 8.450 ;
        RECT 21.785 8.245 21.955 8.450 ;
        RECT 3.465 8.130 3.640 8.245 ;
        RECT 8.045 8.130 8.220 8.245 ;
        RECT 12.625 8.130 12.800 8.245 ;
        RECT 17.205 8.130 17.380 8.245 ;
        RECT 21.785 8.130 21.960 8.245 ;
        RECT 3.470 1.755 3.640 8.130 ;
        RECT 8.050 1.755 8.220 8.130 ;
        RECT 12.630 1.755 12.800 8.130 ;
        RECT 17.210 1.755 17.380 8.130 ;
        RECT 21.790 1.755 21.960 8.130 ;
      LAYER mcon ;
        RECT 3.470 1.835 3.640 8.165 ;
        RECT 8.050 1.835 8.220 8.165 ;
        RECT 12.630 1.835 12.800 8.165 ;
        RECT 17.210 1.835 17.380 8.165 ;
        RECT 21.790 1.835 21.960 8.165 ;
      LAYER met1 ;
        RECT 3.440 1.775 3.670 8.225 ;
        RECT 8.020 1.775 8.250 8.225 ;
        RECT 12.600 1.775 12.830 8.225 ;
        RECT 17.180 1.775 17.410 8.225 ;
        RECT 21.760 1.775 21.990 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 1.180 1.870 1.350 8.245 ;
        RECT 5.760 1.870 5.930 8.245 ;
        RECT 10.340 1.870 10.510 8.245 ;
        RECT 14.920 1.870 15.090 8.245 ;
        RECT 19.500 1.870 19.670 8.245 ;
        RECT 1.175 1.755 1.350 1.870 ;
        RECT 5.755 1.755 5.930 1.870 ;
        RECT 10.335 1.755 10.510 1.870 ;
        RECT 14.915 1.755 15.090 1.870 ;
        RECT 19.495 1.755 19.670 1.870 ;
        RECT 1.175 1.350 1.345 1.755 ;
        RECT 5.755 1.350 5.925 1.755 ;
        RECT 10.335 1.350 10.505 1.755 ;
        RECT 14.915 1.350 15.085 1.755 ;
        RECT 19.495 1.350 19.665 1.755 ;
        RECT 0.940 1.050 22.200 1.350 ;
      LAYER mcon ;
        RECT 1.180 1.835 1.350 8.165 ;
        RECT 5.760 1.835 5.930 8.165 ;
        RECT 10.340 1.835 10.510 8.165 ;
        RECT 14.920 1.835 15.090 8.165 ;
        RECT 19.500 1.835 19.670 8.165 ;
      LAYER met1 ;
        RECT 1.150 1.775 1.380 8.225 ;
        RECT 5.730 1.775 5.960 8.225 ;
        RECT 10.310 1.775 10.540 8.225 ;
        RECT 14.890 1.775 15.120 8.225 ;
        RECT 19.470 1.775 19.700 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 1.470 22.200 9.700 ;
        RECT 0.940 1.465 22.200 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 22.200 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
        RECT 5.840 8.850 6.640 9.250 ;
        RECT 12.340 8.850 13.140 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
        RECT 15.790 9.250 16.090 9.550 ;
        RECT 17.790 9.250 18.090 9.550 ;
        RECT 19.790 9.250 20.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 22.200 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 22.200 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
        RECT 15.790 -0.150 16.090 0.150 ;
        RECT 17.790 -0.150 18.090 0.150 ;
        RECT 19.790 -0.150 20.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 22.200 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9
END LIBRARY

