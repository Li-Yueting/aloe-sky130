magic
tech sky130A
magscale 1 2
timestamp 1654939147
<< pwell >>
rect 120 30 734 1526
<< nmoslvt >>
rect 276 500 676 1500
<< ndiff >>
rect 218 1488 276 1500
rect 218 512 230 1488
rect 264 512 276 1488
rect 218 500 276 512
rect 676 1488 734 1500
rect 676 512 688 1488
rect 722 512 734 1488
rect 676 500 734 512
<< ndiffc >>
rect 230 512 264 1488
rect 688 512 722 1488
<< psubdiff >>
rect 158 160 198 200
rect 158 80 198 120
<< psubdiffcont >>
rect 158 120 198 160
<< poly >>
rect 276 1500 676 1526
rect 276 474 676 500
rect 338 284 458 474
rect 298 264 734 284
rect 298 204 388 264
rect 448 204 734 264
rect 298 184 734 204
<< polycont >>
rect 388 204 448 264
<< locali >>
rect 120 1850 388 1910
rect 448 1850 734 1910
rect 218 1690 734 1750
rect 687 1504 721 1690
rect 230 1488 264 1504
rect 229 512 230 554
rect 687 1488 722 1504
rect 687 1486 688 1488
rect 229 496 264 512
rect 688 496 722 512
rect 229 430 263 496
rect 218 370 734 430
rect 148 160 208 240
rect 298 204 388 264
rect 448 204 734 264
rect 148 120 158 160
rect 198 120 208 160
rect 148 30 208 120
rect 120 -30 388 30
rect 448 -30 734 30
<< viali >>
rect 388 1850 448 1910
rect 230 512 264 1488
rect 688 512 722 1488
rect 388 -30 448 30
<< metal1 >>
rect 120 1910 734 1940
rect 120 1850 388 1910
rect 448 1850 734 1910
rect 120 1820 734 1850
rect 224 1488 270 1500
rect 224 512 230 1488
rect 264 512 270 1488
rect 224 500 270 512
rect 682 1488 728 1500
rect 682 512 688 1488
rect 722 512 728 1488
rect 682 500 728 512
rect 120 30 734 60
rect 120 -30 388 30
rect 448 -30 734 30
rect 120 -60 734 -30
<< labels >>
flabel metal1 218 1850 278 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 218 -30 278 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 674 1690 734 1750 1 FreeSans 800 0 0 0 SOURCE
port 2 n default bidirectional
flabel locali 674 370 734 430 1 FreeSans 800 0 0 0 DRAIN
port 3 n default bidirectional
flabel locali 674 204 734 264 1 FreeSans 800 0 0 0 GATE
port 1 n default bidirectional
<< properties >>
string FIXED_BBOX 0 0 854 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
