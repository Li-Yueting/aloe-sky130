* NGSPICE file created from switch.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136#
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
X0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt transmission_gate en_b out VDD VSS in en
Xsky130_fd_pr__pfet_01v8_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ sky130_fd_pr__pfet_01v8_UNG2NQ
Xsky130_fd_pr__nfet_01v8_6J4AMR_0 out in in out in in VSS out en in out out out sky130_fd_pr__nfet_01v8_6J4AMR
.ends

.subckt sky130_fd_pr__nfet_01v8_E56BNL a_n72_n90# a_16_n90# a_n32_32# VSUBS
X0 a_16_n90# a_n32_32# a_n72_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt switch_5t in en_b VDD out en VSS
Xtransmission_gate_0 en_b transmission_gate_1/in VDD VSS in en transmission_gate
Xtransmission_gate_1 en_b out VDD VSS transmission_gate_1/in en transmission_gate
Xsky130_fd_pr__nfet_01v8_E56BNL_0 VSS transmission_gate_1/in en_b VSS sky130_fd_pr__nfet_01v8_E56BNL
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt my_one_line VDD en in switch_5t_0/en_b en_b out VSS
Xswitch_5t_0 switch_5t_0/in switch_5t_0/en_b VDD out switch_5t_0/en VSS switch_5t
Xtransmission_gate_0 en_b switch_5t_0/in VDD VSS in en transmission_gate
Xsky130_fd_sc_hd__inv_1_0 switch_5t_0/en switch_5t_0/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
.ends

.subckt switch out VSS VDD in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9]
+ in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21]
+ in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] en_b[0] en_b[1]
+ en_b[2] en_b[3] en_b[4] en_b[5] en_b[6] en_b[7] en_b[8] en_b[9] en_b[10] en_b[11]
+ en_b[12] en_b[13] en_b[14] en_b[15] en_b[16] en_b[17] en_b[18] en_b[19] en_b[20]
+ en_b[21] en_b[22] en_b[23] en_b[24] en_b[25] en_b[26] en_b[27] en_b[28] en_b[29]
+ en_b[30] en_b[31] s_en s_en_b
Xmy_one_line_0 VDD s_en in[31] en_b[31] s_en_b out VSS my_one_line
Xmy_one_line_1 VDD s_en in[30] en_b[30] s_en_b out VSS my_one_line
Xmy_one_line_2 VDD s_en in[29] en_b[29] s_en_b out VSS my_one_line
Xmy_one_line_4 VDD s_en in[27] en_b[27] s_en_b out VSS my_one_line
Xmy_one_line_3 VDD s_en in[28] en_b[28] s_en_b out VSS my_one_line
Xmy_one_line_5 VDD s_en in[26] en_b[26] s_en_b out VSS my_one_line
Xmy_one_line_6 VDD s_en in[25] en_b[25] s_en_b out VSS my_one_line
Xmy_one_line_7 VDD s_en in[24] en_b[24] s_en_b out VSS my_one_line
Xmy_one_line_8 VDD s_en in[23] en_b[23] s_en_b out VSS my_one_line
Xmy_one_line_9 VDD s_en in[22] en_b[22] s_en_b out VSS my_one_line
Xmy_one_line_30 VDD s_en in[1] en_b[1] s_en_b out VSS my_one_line
Xmy_one_line_31 VDD s_en in[0] en_b[0] s_en_b out VSS my_one_line
Xmy_one_line_20 VDD s_en in[11] en_b[11] s_en_b out VSS my_one_line
Xmy_one_line_22 VDD s_en in[9] en_b[9] s_en_b out VSS my_one_line
Xmy_one_line_21 VDD s_en in[10] en_b[10] s_en_b out VSS my_one_line
Xmy_one_line_11 VDD s_en in[20] en_b[20] s_en_b out VSS my_one_line
Xmy_one_line_10 VDD s_en in[21] en_b[21] s_en_b out VSS my_one_line
Xmy_one_line_23 VDD s_en in[8] en_b[8] s_en_b out VSS my_one_line
Xmy_one_line_12 VDD s_en in[19] en_b[19] s_en_b out VSS my_one_line
Xmy_one_line_24 VDD s_en in[7] en_b[7] s_en_b out VSS my_one_line
Xmy_one_line_13 VDD s_en in[18] en_b[18] s_en_b out VSS my_one_line
Xmy_one_line_25 VDD s_en in[6] en_b[6] s_en_b out VSS my_one_line
Xmy_one_line_14 VDD s_en in[17] en_b[17] s_en_b out VSS my_one_line
Xmy_one_line_26 VDD s_en in[5] en_b[5] s_en_b out VSS my_one_line
Xmy_one_line_15 VDD s_en in[16] en_b[16] s_en_b out VSS my_one_line
Xmy_one_line_27 VDD s_en in[4] en_b[4] s_en_b out VSS my_one_line
Xmy_one_line_16 VDD s_en in[15] en_b[15] s_en_b out VSS my_one_line
Xmy_one_line_28 VDD s_en in[3] en_b[3] s_en_b out VSS my_one_line
Xmy_one_line_17 VDD s_en in[14] en_b[14] s_en_b out VSS my_one_line
Xmy_one_line_29 VDD s_en in[2] en_b[2] s_en_b out VSS my_one_line
Xmy_one_line_19 VDD s_en in[12] en_b[12] s_en_b out VSS my_one_line
Xmy_one_line_18 VDD s_en in[13] en_b[13] s_en_b out VSS my_one_line
.ends

