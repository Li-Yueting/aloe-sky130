VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_7
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_7 ;
  ORIGIN 0.000 0.000 ;
  SIZE 46.900 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 80.919998 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.965 5.085 6.435 ;
        RECT 8.315 2.965 11.785 6.435 ;
        RECT 15.015 2.965 18.485 6.435 ;
        RECT 21.715 2.965 25.185 6.435 ;
        RECT 28.415 2.965 31.885 6.435 ;
        RECT 35.115 2.965 38.585 6.435 ;
        RECT 41.815 2.965 45.285 6.435 ;
      LAYER mcon ;
        RECT 1.980 5.830 2.150 6.000 ;
        RECT 2.480 5.830 2.650 6.000 ;
        RECT 2.980 5.830 3.150 6.000 ;
        RECT 3.480 5.830 3.650 6.000 ;
        RECT 3.980 5.830 4.150 6.000 ;
        RECT 4.480 5.830 4.650 6.000 ;
        RECT 1.980 5.330 2.150 5.500 ;
        RECT 2.480 5.330 2.650 5.500 ;
        RECT 2.980 5.330 3.150 5.500 ;
        RECT 3.480 5.330 3.650 5.500 ;
        RECT 3.980 5.330 4.150 5.500 ;
        RECT 4.480 5.330 4.650 5.500 ;
        RECT 1.980 4.830 2.150 5.000 ;
        RECT 2.480 4.830 2.650 5.000 ;
        RECT 2.980 4.830 3.150 5.000 ;
        RECT 3.480 4.830 3.650 5.000 ;
        RECT 3.980 4.830 4.150 5.000 ;
        RECT 4.480 4.830 4.650 5.000 ;
        RECT 1.980 4.330 2.150 4.500 ;
        RECT 2.480 4.330 2.650 4.500 ;
        RECT 2.980 4.330 3.150 4.500 ;
        RECT 3.480 4.330 3.650 4.500 ;
        RECT 3.980 4.330 4.150 4.500 ;
        RECT 4.480 4.330 4.650 4.500 ;
        RECT 1.980 3.830 2.150 4.000 ;
        RECT 2.480 3.830 2.650 4.000 ;
        RECT 2.980 3.830 3.150 4.000 ;
        RECT 3.480 3.830 3.650 4.000 ;
        RECT 3.980 3.830 4.150 4.000 ;
        RECT 4.480 3.830 4.650 4.000 ;
        RECT 1.980 3.330 2.150 3.500 ;
        RECT 2.480 3.330 2.650 3.500 ;
        RECT 2.980 3.330 3.150 3.500 ;
        RECT 3.480 3.330 3.650 3.500 ;
        RECT 3.980 3.330 4.150 3.500 ;
        RECT 4.480 3.330 4.650 3.500 ;
        RECT 8.680 5.830 8.850 6.000 ;
        RECT 9.180 5.830 9.350 6.000 ;
        RECT 9.680 5.830 9.850 6.000 ;
        RECT 10.180 5.830 10.350 6.000 ;
        RECT 10.680 5.830 10.850 6.000 ;
        RECT 11.180 5.830 11.350 6.000 ;
        RECT 8.680 5.330 8.850 5.500 ;
        RECT 9.180 5.330 9.350 5.500 ;
        RECT 9.680 5.330 9.850 5.500 ;
        RECT 10.180 5.330 10.350 5.500 ;
        RECT 10.680 5.330 10.850 5.500 ;
        RECT 11.180 5.330 11.350 5.500 ;
        RECT 8.680 4.830 8.850 5.000 ;
        RECT 9.180 4.830 9.350 5.000 ;
        RECT 9.680 4.830 9.850 5.000 ;
        RECT 10.180 4.830 10.350 5.000 ;
        RECT 10.680 4.830 10.850 5.000 ;
        RECT 11.180 4.830 11.350 5.000 ;
        RECT 8.680 4.330 8.850 4.500 ;
        RECT 9.180 4.330 9.350 4.500 ;
        RECT 9.680 4.330 9.850 4.500 ;
        RECT 10.180 4.330 10.350 4.500 ;
        RECT 10.680 4.330 10.850 4.500 ;
        RECT 11.180 4.330 11.350 4.500 ;
        RECT 8.680 3.830 8.850 4.000 ;
        RECT 9.180 3.830 9.350 4.000 ;
        RECT 9.680 3.830 9.850 4.000 ;
        RECT 10.180 3.830 10.350 4.000 ;
        RECT 10.680 3.830 10.850 4.000 ;
        RECT 11.180 3.830 11.350 4.000 ;
        RECT 8.680 3.330 8.850 3.500 ;
        RECT 9.180 3.330 9.350 3.500 ;
        RECT 9.680 3.330 9.850 3.500 ;
        RECT 10.180 3.330 10.350 3.500 ;
        RECT 10.680 3.330 10.850 3.500 ;
        RECT 11.180 3.330 11.350 3.500 ;
        RECT 15.380 5.830 15.550 6.000 ;
        RECT 15.880 5.830 16.050 6.000 ;
        RECT 16.380 5.830 16.550 6.000 ;
        RECT 16.880 5.830 17.050 6.000 ;
        RECT 17.380 5.830 17.550 6.000 ;
        RECT 17.880 5.830 18.050 6.000 ;
        RECT 15.380 5.330 15.550 5.500 ;
        RECT 15.880 5.330 16.050 5.500 ;
        RECT 16.380 5.330 16.550 5.500 ;
        RECT 16.880 5.330 17.050 5.500 ;
        RECT 17.380 5.330 17.550 5.500 ;
        RECT 17.880 5.330 18.050 5.500 ;
        RECT 15.380 4.830 15.550 5.000 ;
        RECT 15.880 4.830 16.050 5.000 ;
        RECT 16.380 4.830 16.550 5.000 ;
        RECT 16.880 4.830 17.050 5.000 ;
        RECT 17.380 4.830 17.550 5.000 ;
        RECT 17.880 4.830 18.050 5.000 ;
        RECT 15.380 4.330 15.550 4.500 ;
        RECT 15.880 4.330 16.050 4.500 ;
        RECT 16.380 4.330 16.550 4.500 ;
        RECT 16.880 4.330 17.050 4.500 ;
        RECT 17.380 4.330 17.550 4.500 ;
        RECT 17.880 4.330 18.050 4.500 ;
        RECT 15.380 3.830 15.550 4.000 ;
        RECT 15.880 3.830 16.050 4.000 ;
        RECT 16.380 3.830 16.550 4.000 ;
        RECT 16.880 3.830 17.050 4.000 ;
        RECT 17.380 3.830 17.550 4.000 ;
        RECT 17.880 3.830 18.050 4.000 ;
        RECT 15.380 3.330 15.550 3.500 ;
        RECT 15.880 3.330 16.050 3.500 ;
        RECT 16.380 3.330 16.550 3.500 ;
        RECT 16.880 3.330 17.050 3.500 ;
        RECT 17.380 3.330 17.550 3.500 ;
        RECT 17.880 3.330 18.050 3.500 ;
        RECT 22.080 5.830 22.250 6.000 ;
        RECT 22.580 5.830 22.750 6.000 ;
        RECT 23.080 5.830 23.250 6.000 ;
        RECT 23.580 5.830 23.750 6.000 ;
        RECT 24.080 5.830 24.250 6.000 ;
        RECT 24.580 5.830 24.750 6.000 ;
        RECT 22.080 5.330 22.250 5.500 ;
        RECT 22.580 5.330 22.750 5.500 ;
        RECT 23.080 5.330 23.250 5.500 ;
        RECT 23.580 5.330 23.750 5.500 ;
        RECT 24.080 5.330 24.250 5.500 ;
        RECT 24.580 5.330 24.750 5.500 ;
        RECT 22.080 4.830 22.250 5.000 ;
        RECT 22.580 4.830 22.750 5.000 ;
        RECT 23.080 4.830 23.250 5.000 ;
        RECT 23.580 4.830 23.750 5.000 ;
        RECT 24.080 4.830 24.250 5.000 ;
        RECT 24.580 4.830 24.750 5.000 ;
        RECT 22.080 4.330 22.250 4.500 ;
        RECT 22.580 4.330 22.750 4.500 ;
        RECT 23.080 4.330 23.250 4.500 ;
        RECT 23.580 4.330 23.750 4.500 ;
        RECT 24.080 4.330 24.250 4.500 ;
        RECT 24.580 4.330 24.750 4.500 ;
        RECT 22.080 3.830 22.250 4.000 ;
        RECT 22.580 3.830 22.750 4.000 ;
        RECT 23.080 3.830 23.250 4.000 ;
        RECT 23.580 3.830 23.750 4.000 ;
        RECT 24.080 3.830 24.250 4.000 ;
        RECT 24.580 3.830 24.750 4.000 ;
        RECT 22.080 3.330 22.250 3.500 ;
        RECT 22.580 3.330 22.750 3.500 ;
        RECT 23.080 3.330 23.250 3.500 ;
        RECT 23.580 3.330 23.750 3.500 ;
        RECT 24.080 3.330 24.250 3.500 ;
        RECT 24.580 3.330 24.750 3.500 ;
        RECT 28.780 5.830 28.950 6.000 ;
        RECT 29.280 5.830 29.450 6.000 ;
        RECT 29.780 5.830 29.950 6.000 ;
        RECT 30.280 5.830 30.450 6.000 ;
        RECT 30.780 5.830 30.950 6.000 ;
        RECT 31.280 5.830 31.450 6.000 ;
        RECT 28.780 5.330 28.950 5.500 ;
        RECT 29.280 5.330 29.450 5.500 ;
        RECT 29.780 5.330 29.950 5.500 ;
        RECT 30.280 5.330 30.450 5.500 ;
        RECT 30.780 5.330 30.950 5.500 ;
        RECT 31.280 5.330 31.450 5.500 ;
        RECT 28.780 4.830 28.950 5.000 ;
        RECT 29.280 4.830 29.450 5.000 ;
        RECT 29.780 4.830 29.950 5.000 ;
        RECT 30.280 4.830 30.450 5.000 ;
        RECT 30.780 4.830 30.950 5.000 ;
        RECT 31.280 4.830 31.450 5.000 ;
        RECT 28.780 4.330 28.950 4.500 ;
        RECT 29.280 4.330 29.450 4.500 ;
        RECT 29.780 4.330 29.950 4.500 ;
        RECT 30.280 4.330 30.450 4.500 ;
        RECT 30.780 4.330 30.950 4.500 ;
        RECT 31.280 4.330 31.450 4.500 ;
        RECT 28.780 3.830 28.950 4.000 ;
        RECT 29.280 3.830 29.450 4.000 ;
        RECT 29.780 3.830 29.950 4.000 ;
        RECT 30.280 3.830 30.450 4.000 ;
        RECT 30.780 3.830 30.950 4.000 ;
        RECT 31.280 3.830 31.450 4.000 ;
        RECT 28.780 3.330 28.950 3.500 ;
        RECT 29.280 3.330 29.450 3.500 ;
        RECT 29.780 3.330 29.950 3.500 ;
        RECT 30.280 3.330 30.450 3.500 ;
        RECT 30.780 3.330 30.950 3.500 ;
        RECT 31.280 3.330 31.450 3.500 ;
        RECT 35.480 5.830 35.650 6.000 ;
        RECT 35.980 5.830 36.150 6.000 ;
        RECT 36.480 5.830 36.650 6.000 ;
        RECT 36.980 5.830 37.150 6.000 ;
        RECT 37.480 5.830 37.650 6.000 ;
        RECT 37.980 5.830 38.150 6.000 ;
        RECT 35.480 5.330 35.650 5.500 ;
        RECT 35.980 5.330 36.150 5.500 ;
        RECT 36.480 5.330 36.650 5.500 ;
        RECT 36.980 5.330 37.150 5.500 ;
        RECT 37.480 5.330 37.650 5.500 ;
        RECT 37.980 5.330 38.150 5.500 ;
        RECT 35.480 4.830 35.650 5.000 ;
        RECT 35.980 4.830 36.150 5.000 ;
        RECT 36.480 4.830 36.650 5.000 ;
        RECT 36.980 4.830 37.150 5.000 ;
        RECT 37.480 4.830 37.650 5.000 ;
        RECT 37.980 4.830 38.150 5.000 ;
        RECT 35.480 4.330 35.650 4.500 ;
        RECT 35.980 4.330 36.150 4.500 ;
        RECT 36.480 4.330 36.650 4.500 ;
        RECT 36.980 4.330 37.150 4.500 ;
        RECT 37.480 4.330 37.650 4.500 ;
        RECT 37.980 4.330 38.150 4.500 ;
        RECT 35.480 3.830 35.650 4.000 ;
        RECT 35.980 3.830 36.150 4.000 ;
        RECT 36.480 3.830 36.650 4.000 ;
        RECT 36.980 3.830 37.150 4.000 ;
        RECT 37.480 3.830 37.650 4.000 ;
        RECT 37.980 3.830 38.150 4.000 ;
        RECT 35.480 3.330 35.650 3.500 ;
        RECT 35.980 3.330 36.150 3.500 ;
        RECT 36.480 3.330 36.650 3.500 ;
        RECT 36.980 3.330 37.150 3.500 ;
        RECT 37.480 3.330 37.650 3.500 ;
        RECT 37.980 3.330 38.150 3.500 ;
        RECT 42.180 5.830 42.350 6.000 ;
        RECT 42.680 5.830 42.850 6.000 ;
        RECT 43.180 5.830 43.350 6.000 ;
        RECT 43.680 5.830 43.850 6.000 ;
        RECT 44.180 5.830 44.350 6.000 ;
        RECT 44.680 5.830 44.850 6.000 ;
        RECT 42.180 5.330 42.350 5.500 ;
        RECT 42.680 5.330 42.850 5.500 ;
        RECT 43.180 5.330 43.350 5.500 ;
        RECT 43.680 5.330 43.850 5.500 ;
        RECT 44.180 5.330 44.350 5.500 ;
        RECT 44.680 5.330 44.850 5.500 ;
        RECT 42.180 4.830 42.350 5.000 ;
        RECT 42.680 4.830 42.850 5.000 ;
        RECT 43.180 4.830 43.350 5.000 ;
        RECT 43.680 4.830 43.850 5.000 ;
        RECT 44.180 4.830 44.350 5.000 ;
        RECT 44.680 4.830 44.850 5.000 ;
        RECT 42.180 4.330 42.350 4.500 ;
        RECT 42.680 4.330 42.850 4.500 ;
        RECT 43.180 4.330 43.350 4.500 ;
        RECT 43.680 4.330 43.850 4.500 ;
        RECT 44.180 4.330 44.350 4.500 ;
        RECT 44.680 4.330 44.850 4.500 ;
        RECT 42.180 3.830 42.350 4.000 ;
        RECT 42.680 3.830 42.850 4.000 ;
        RECT 43.180 3.830 43.350 4.000 ;
        RECT 43.680 3.830 43.850 4.000 ;
        RECT 44.180 3.830 44.350 4.000 ;
        RECT 44.680 3.830 44.850 4.000 ;
        RECT 42.180 3.330 42.350 3.500 ;
        RECT 42.680 3.330 42.850 3.500 ;
        RECT 43.180 3.330 43.350 3.500 ;
        RECT 43.680 3.330 43.850 3.500 ;
        RECT 44.180 3.330 44.350 3.500 ;
        RECT 44.680 3.330 44.850 3.500 ;
      LAYER met1 ;
        RECT 1.820 3.170 45.310 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 187.102295 ;
    ANTENNADIFFAREA 138.823303 ;
    PORT
      LAYER pwell ;
        RECT 0.000 7.285 46.900 8.050 ;
        RECT 0.000 2.115 0.765 7.285 ;
        RECT 5.935 2.115 7.465 7.285 ;
        RECT 12.635 2.115 14.165 7.285 ;
        RECT 19.335 2.115 20.865 7.285 ;
        RECT 26.035 2.115 27.565 7.285 ;
        RECT 32.735 2.115 34.265 7.285 ;
        RECT 39.435 2.115 40.965 7.285 ;
        RECT 46.135 2.115 46.900 7.285 ;
        RECT 0.000 1.350 46.900 2.115 ;
      LAYER li1 ;
        RECT 0.130 7.050 46.785 7.920 ;
        RECT 0.130 2.350 0.625 7.050 ;
        RECT 0.945 6.745 5.755 7.050 ;
        RECT 0.945 2.655 1.305 6.745 ;
        RECT 5.395 2.655 5.755 6.745 ;
        RECT 0.945 2.350 5.755 2.655 ;
        RECT 6.075 2.350 7.325 7.050 ;
        RECT 7.645 6.745 12.455 7.050 ;
        RECT 7.645 2.655 8.005 6.745 ;
        RECT 12.095 2.655 12.455 6.745 ;
        RECT 7.645 2.350 12.455 2.655 ;
        RECT 12.775 2.350 14.025 7.050 ;
        RECT 14.345 6.745 19.155 7.050 ;
        RECT 14.345 2.655 14.705 6.745 ;
        RECT 18.795 2.655 19.155 6.745 ;
        RECT 14.345 2.350 19.155 2.655 ;
        RECT 19.475 2.350 20.725 7.050 ;
        RECT 21.045 6.745 25.855 7.050 ;
        RECT 21.045 2.655 21.405 6.745 ;
        RECT 25.495 2.655 25.855 6.745 ;
        RECT 21.045 2.350 25.855 2.655 ;
        RECT 26.175 2.350 27.425 7.050 ;
        RECT 27.745 6.745 32.555 7.050 ;
        RECT 27.745 2.655 28.105 6.745 ;
        RECT 32.195 2.655 32.555 6.745 ;
        RECT 27.745 2.350 32.555 2.655 ;
        RECT 32.875 2.350 34.125 7.050 ;
        RECT 34.445 6.745 39.255 7.050 ;
        RECT 34.445 2.655 34.805 6.745 ;
        RECT 38.895 2.655 39.255 6.745 ;
        RECT 34.445 2.350 39.255 2.655 ;
        RECT 39.575 2.350 40.825 7.050 ;
        RECT 41.145 6.745 45.955 7.050 ;
        RECT 41.145 2.655 41.505 6.745 ;
        RECT 45.595 2.655 45.955 6.745 ;
        RECT 41.145 2.350 45.955 2.655 ;
        RECT 46.275 2.350 46.770 7.050 ;
        RECT 0.130 1.480 46.785 2.350 ;
    END
  END Base
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 46.900 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 1.850 9.250 2.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 3.850 9.250 4.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 5.850 9.250 6.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 7.850 9.250 8.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 9.850 9.250 10.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 11.850 9.250 12.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 13.850 9.250 14.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 15.850 9.250 16.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 17.850 9.250 18.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
        RECT 19.850 9.250 20.150 9.550 ;
        RECT 20.850 9.250 21.150 9.550 ;
        RECT 21.850 9.250 22.150 9.550 ;
        RECT 22.850 9.250 23.150 9.550 ;
        RECT 23.850 9.250 24.150 9.550 ;
        RECT 24.850 9.250 25.150 9.550 ;
        RECT 25.850 9.250 26.150 9.550 ;
        RECT 26.850 9.250 27.150 9.550 ;
        RECT 27.850 9.250 28.150 9.550 ;
        RECT 28.850 9.250 29.150 9.550 ;
        RECT 29.850 9.250 30.150 9.550 ;
        RECT 30.850 9.250 31.150 9.550 ;
        RECT 31.850 9.250 32.150 9.550 ;
        RECT 32.850 9.250 33.150 9.550 ;
        RECT 33.850 9.250 34.150 9.550 ;
        RECT 34.850 9.250 35.150 9.550 ;
        RECT 35.850 9.250 36.150 9.550 ;
        RECT 36.850 9.250 37.150 9.550 ;
        RECT 37.850 9.250 38.150 9.550 ;
        RECT 38.850 9.250 39.150 9.550 ;
        RECT 39.850 9.250 40.150 9.550 ;
        RECT 40.850 9.250 41.150 9.550 ;
        RECT 41.850 9.250 42.150 9.550 ;
        RECT 42.850 9.250 43.150 9.550 ;
        RECT 43.850 9.250 44.150 9.550 ;
        RECT 44.850 9.250 45.150 9.550 ;
        RECT 45.850 9.250 46.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 46.900 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 46.900 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.850 -0.150 21.150 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.850 -0.150 23.150 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.850 -0.150 25.150 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.850 -0.150 27.150 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.850 -0.150 29.150 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.850 -0.150 31.150 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.850 -0.150 33.150 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.850 -0.150 35.150 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.850 -0.150 37.150 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.850 -0.150 39.150 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.850 -0.150 41.150 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.850 -0.150 43.150 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.850 -0.150 45.150 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 46.900 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_7
END LIBRARY

