magic
tech sky130A
magscale 1 2
timestamp 1651598395
<< nwell >>
rect 0 293 588 1940
<< pmoslvt >>
rect 94 355 494 1645
<< pdiff >>
rect 36 1633 94 1645
rect 36 367 48 1633
rect 82 367 94 1633
rect 36 355 94 367
rect 494 1633 552 1645
rect 494 367 506 1633
rect 540 367 552 1633
rect 494 355 552 367
<< pdiffc >>
rect 48 367 82 1633
rect 506 367 540 1633
<< poly >>
rect 94 1645 494 1671
rect 94 329 494 355
rect 240 184 360 329
rect 0 164 588 184
rect 0 104 170 164
rect 230 104 588 164
rect 0 84 588 104
<< polycont >>
rect 170 104 230 164
<< locali >>
rect 0 1850 170 1910
rect 230 1850 588 1910
rect 0 1730 588 1790
rect 505 1649 539 1730
rect 48 1633 82 1649
rect 47 367 48 374
rect 505 1633 540 1649
rect 505 1626 506 1633
rect 47 351 82 367
rect 506 351 540 367
rect 47 270 81 351
rect 0 210 588 270
rect 0 104 170 164
rect 230 104 588 164
rect 0 -30 170 30
rect 230 -30 588 30
<< viali >>
rect 170 1850 230 1910
rect 48 367 82 1633
rect 506 367 540 1633
rect 170 -30 230 30
<< metal1 >>
rect 0 1910 588 1940
rect 0 1850 170 1910
rect 230 1850 588 1910
rect 0 1820 588 1850
rect 42 1633 88 1645
rect 42 367 48 1633
rect 82 367 88 1633
rect 42 355 88 367
rect 500 1633 546 1645
rect 500 367 506 1633
rect 540 367 546 1633
rect 500 355 546 367
rect 0 30 588 60
rect 0 -30 170 30
rect 230 -30 588 30
rect 0 -60 588 -30
<< labels >>
flabel nwell 170 1850 230 1910 1 FreeSans 800 0 0 0 VPB
port 4 n power bidirectional
flabel metal1 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 5 n power bidirectional
flabel metal1 0 -30 60 30 1 FreeSans 800 0 0 0 VGND
port 6 n ground bidirectional
flabel locali 528 1730 588 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 528 210 588 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 528 104 588 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 588 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
