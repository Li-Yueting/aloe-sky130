
* NGSPICE file created from bgr_top.ext - technology: sky130A

.subckt sky130_asc_res_xhigh_po_2p85_1 Rin Rout VPWR VGND a_2148_115#
X0 Rin a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X1 Rout a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
C0 Rin VPWR 0.17fF
C1 Rout Rin 0.12fF
C2 a_2148_115# VPWR 0.17fF
C3 VPWR VGND 2.31fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2148_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_60 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.79855e+13p pd=4.1788e+08u as=5.6115e+13p ps=4.044e+08u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X12 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X13 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X14 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X15 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X16 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X17 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X18 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X19 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X20 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X21 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X22 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X23 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X24 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X26 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X27 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X28 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X29 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X30 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X31 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X32 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X33 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X34 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X35 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X36 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X37 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X38 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X39 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X40 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X41 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X42 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X43 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X44 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X45 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X46 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X47 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X48 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X50 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X51 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X52 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X53 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X54 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X55 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X56 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X58 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X59 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 VPWR SOURCE 22.83fF
C1 VGND SOURCE 0.32fF
C2 GATE SOURCE 0.18fF
C3 DRAIN SOURCE 1.25fF
C4 GATE VPWR 27.32fF
C5 GATE VGND 12.31fF
C6 DRAIN VPWR 1.83fF
C7 DRAIN VGND 5.28fF
C8 DRAIN GATE 25.46fF
C9 VGND VSUBS 25.41fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 9.62fF
C12 GATE VSUBS 30.27fF
C13 VPWR VSUBS 142.65fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_7 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
C0 Base Emitter 18.67fF
C1 VGND Collector 9.81fF
C2 VPWR Collector 11.49fF
C3 Emitter Collector 9.06fF
C4 Base Collector 28.86fF
.ends

.subckt sky130_asc_res_xhigh_po_2p85_2 Rin Rout VPWR a_2723_115# VGND
X0 Rout a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X1 Rin a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
C0 Rin Rout 0.12fF
C1 VPWR Rin 0.17fF
C2 a_2723_115# VPWR 0.17fF
C3 VPWR VGND 2.83fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2723_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_12 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=1.1223e+13p pd=8.088e+07u as=1.30935e+13p ps=9.436e+07u w=6.45e+06u l=2e+06u
X1 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 VPWR DRAIN 0.42fF
C1 GATE DRAIN 5.17fF
C2 GATE VPWR 5.46fF
C3 VGND DRAIN 1.08fF
C4 SOURCE DRAIN 0.26fF
C5 SOURCE VPWR 4.54fF
C6 VGND GATE 2.51fF
C7 SOURCE GATE 0.04fF
C8 SOURCE VGND 0.06fF
C9 VGND VSUBS 5.31fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.99fF
C12 GATE VSUBS 6.20fF
C13 VPWR VSUBS 29.52fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_9 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=5.8e+12p pd=4.29e+07u as=5.8e+12p ps=4.29e+07u w=4e+06u l=2e+06u
X1 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
C0 SOURCE GATE 0.01fF
C1 DRAIN GATE 1.66fF
C2 DRAIN SOURCE 0.05fF
C3 VPWR SOURCE 1.38fF
C4 VPWR VGND 3.99fF
C5 SOURCE VGND 2.64fF
C6 DRAIN VGND 2.28fF
C7 GATE VGND 11.48fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_6 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.6115e+12p pd=4.044e+07u as=7.482e+12p ps=5.392e+07u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 DRAIN VGND 0.56fF
C1 SOURCE VGND 0.03fF
C2 SOURCE DRAIN 0.14fF
C3 GATE VGND 1.28fF
C4 GATE DRAIN 2.63fF
C5 VPWR DRAIN 0.24fF
C6 GATE SOURCE 0.02fF
C7 VPWR SOURCE 2.27fF
C8 VPWR GATE 2.73fF
C9 VGND VSUBS 2.79fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.04fF
C12 GATE VSUBS 3.19fF
C13 VPWR VSUBS 15.38fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_1 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
C0 Emitter Base 1.55fF
C1 VGND Collector 1.50fF
C2 VPWR Collector 1.46fF
C3 Emitter Collector 0.40fF
C4 Base Collector 3.33fF
.ends

.subckt sky130_asc_cap_mim_m3_1 Cin Cout VPWR VGND VSUBS
X0 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X9 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X10 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X13 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X15 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
C0 Cout Cin 28.31fF
C1 Cout VSUBS 2.81fF
C2 Cin VSUBS 6.38fF
C3 VGND VSUBS 6.63fF
C4 VPWR VSUBS 6.63fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_8 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X7 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
C0 Base Emitter 21.50fF
C1 VGND Collector 11.20fF
C2 VPWR Collector 13.12fF
C3 Emitter Collector 10.49fF
C4 Base Collector 33.06fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
C0 GATE SOURCE 0.00fF
C1 SOURCE DRAIN 0.01fF
C2 VPWR SOURCE 0.17fF
C3 GATE DRAIN 0.18fF
C4 VPWR VGND 0.64fF
C5 SOURCE VGND 0.40fF
C6 DRAIN VGND 0.34fF
C7 GATE VGND 1.34fF
.ends

.subckt bgr_top porst va vb vbg VSS VDD
Xsky130_asc_res_xhigh_po_2p85_1_7 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_8 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_9 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_60_0 sky130_asc_cap_mim_m3_1_4/Cout VDD vbg VSS VDD VSS
+ sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_1 sky130_asc_cap_mim_m3_1_4/Cout VDD vb VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_2 sky130_asc_cap_mim_m3_1_4/Cout VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_res_xhigh_po_2p85_1_30 va sky130_asc_res_xhigh_po_2p85_1_29/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_20 vb sky130_asc_res_xhigh_po_2p85_1_19/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_7_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_7
Xsky130_asc_res_xhigh_po_2p85_1_10 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_21 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_0 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_11 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_1 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_12 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_23 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_13 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_0 VDD VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_25 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_14 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_1 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_26 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_15 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_16 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_27 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_17 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_28 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_0 porst VSS sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_18 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_29 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_0 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_cap_mim_m3_1_4/Cout
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_nfet_01v8_lvt_9_1 va sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_cap_mim_m3_1_4/Cout
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_19 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_1 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_pnp_05v5_W3p40L3p40_1_0 va VSS VSS VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_1
Xsky130_asc_nfet_01v8_lvt_9_2 vb sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_cap_mim_m3_1_0 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_1 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_2 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_1 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_3 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_2 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_4 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_3 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_5 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_0 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_6 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_0 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_1 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_7 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_1 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_2 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_8 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_3 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_9 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_4 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_5 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_6 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
X0 sky130_asc_pfet_01v8_lvt_6_1/GATE.t1 sky130_asc_pfet_01v8_lvt_6_1/GATE.t0 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.02014e+14p ps=1.45584e+09u w=0u l=0u
X1 sky130_asc_nfet_01v8_lvt_1_1/DRAIN va.t7 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=1.276e+13p pd=9.438e+07u as=1.16e+13p ps=8.58e+07u w=0u l=0u
X2 VSS.t186 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X3 va VDD.t12 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=8.2639e+13p pd=5.2584e+08u as=0p ps=0u w=0u l=0u
X4 VSS VSS.t26 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X5 VSS VSS.t34 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X6 VSS.t191 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X7 VSS.t150 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X8 va VDD.t0 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X9 VSS.t134 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X10 VSS.t135 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X11 VSS.t217 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X12 VSS.t141 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X13 VSS VSS.t66 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X14 VSS.t177 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X15 VSS.t219 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X16 VSS.t174 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X17 VSS.t184 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X18 sky130_asc_pfet_01v8_lvt_6_1/GATE.t5 sky130_asc_pfet_01v8_lvt_6_1/GATE.t4 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X19 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE.t2 sky130_asc_pfet_01v8_lvt_6_1/GATE.t3 VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 VSS VSS.t6 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X21 VSS.t179 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X22 VSS VSS.t62 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X23 VSS.t195 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X24 VSS.t144 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X25 VSS.t203 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X26 VSS.t133 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X27 VDD.t5 VDD.t3 va VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X28 va VDD.t9 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X29 VSS VSS.t48 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X30 VSS.t204 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X31 VSS VSS.t64 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X32 VSS VSS.t46 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X33 VSS VSS.t10 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X34 va VDD.t27 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X35 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE.t10 sky130_asc_pfet_01v8_lvt_6_1/GATE.t11 VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X36 VSS.t192 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X37 VSS.t173 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X38 VSS.t149 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X39 VSS VSS.t18 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X40 sky130_asc_cap_mim_m3_1_4/Cout porst.t2 VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.6444e+14p ps=1.48406e+09u w=0u l=0u
X41 VSS VSS.t32 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X42 VDD.t35 VDD.t33 va VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X43 VSS porst.t7 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X44 VSS.t193 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X45 VSS VSS.t76 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X46 VSS.t138 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X47 VSS.t212 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X48 VDD.t17 VDD.t15 va VDD.t16 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X49 VSS.t136 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X50 VSS VSS.t60 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X51 VSS.t129 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X52 VSS.t178 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X53 VSS porst.t5 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X54 VSS.t122 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X55 VSS.t183 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X56 VSS.t176 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X57 VSS.t190 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X58 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE.t8 sky130_asc_pfet_01v8_lvt_6_1/GATE.t9 VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X59 VSS.t208 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X60 VSS VSS.t44 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X61 VSS.t168 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X62 VSS VSS.t68 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X63 VSS VSS.t52 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X64 VSS VSS.t30 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X65 VSS.t205 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X66 VSS.t182 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X67 VSS.t127 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X68 VSS.t140 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X69 VSS.t153 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X70 VSS VSS.t2 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X71 VSS.t210 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X72 VSS VSS.t74 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X73 VSS VSS.t56 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X74 VSS VSS.t16 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X75 VSS.t120 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X76 VSS.t167 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X77 VSS VSS.t36 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X78 VSS porst.t1 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X79 sky130_asc_cap_mim_m3_1_4/Cout porst.t8 VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X80 VSS.t148 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X81 VSS.t201 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X82 VSS.t161 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X83 VSS porst.t3 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X84 sky130_asc_cap_mim_m3_1_4/Cout porst.t6 VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X85 VSS.t180 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X86 VSS VSS.t40 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X87 VSS.t155 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X88 VSS.t181 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X89 VSS.t143 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X90 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE.t16 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=7.482e+12p ps=5.392e+07u w=0u l=0u
X91 VSS.t137 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X92 VSS.t151 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X93 VSS porst.t0 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X94 VSS VSS.t28 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X95 VSS.t206 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X96 VSS VSS.t14 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X97 VSS.t157 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X98 VSS.t139 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X99 sky130_asc_nfet_01v8_lvt_1_1/DRAIN vb.t1 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+12p ps=4.29e+07u w=0u l=0u
X100 VSS.t185 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X101 sky130_asc_nfet_01v8_lvt_1_1/DRAIN va.t3 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X102 VSS.t211 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X103 VSS.t166 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X104 VSS.t171 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X105 sky130_asc_pfet_01v8_lvt_6_1/GATE vb.t2 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X106 sky130_asc_nfet_01v8_lvt_1_1/DRAIN vb.t3 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X107 VSS VSS.t0 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X108 VSS.t123 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X109 VSS.t194 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X110 VSS.t189 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X111 VSS.t199 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X112 VSS VSS.t20 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X113 VSS.t124 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X114 VSS.t214 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X115 VSS.t163 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X116 sky130_asc_cap_mim_m3_1_4/Cout porst.t4 VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X117 VSS VSS.t24 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X118 VSS.t215 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X119 VSS.t146 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X120 sky130_asc_nfet_01v8_lvt_1_1/DRAIN vb.t5 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X121 VSS.t164 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X122 VSS.t152 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X123 VSS.t175 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X124 sky130_asc_cap_mim_m3_1_4/Cout va.t2 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X125 sky130_asc_nfet_01v8_lvt_1_1/DRAIN vb.t7 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X126 VSS VSS.t12 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X127 VSS.t132 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X128 VSS.t154 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X129 VSS VSS.t54 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X130 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE.t13 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X131 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_pfet_01v8_lvt_6_1/GATE.t17 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X132 VSS.t213 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X133 sky130_asc_cap_mim_m3_1_4/Cout va.t4 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X134 sky130_asc_nfet_01v8_lvt_1_1/DRAIN va.t5 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X135 VSS.t172 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X136 va VDD.t30 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X137 VDD.t26 VDD.t24 va VDD.t25 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X138 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_pfet_01v8_lvt_6_1/GATE.t15 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X139 VSS.t147 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X140 VSS.t198 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X141 VSS.t159 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X142 sky130_asc_cap_mim_m3_1_4/Cout va.t8 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X143 VSS VSS.t78 va sky130_fd_pr__pnp_05v5 area=0p
X144 sky130_asc_pfet_01v8_lvt_6_1/GATE vb.t8 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X145 VSS VSS.t38 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X146 VSS VSS.t4 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X147 VSS.t128 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X148 sky130_asc_nfet_01v8_lvt_1_1/DRAIN va.t1 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X149 VSS VSS.t58 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X150 VSS.t196 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X151 VSS VSS.t72 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X152 sky130_asc_pfet_01v8_lvt_6_1/GATE vb.t6 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X153 VSS.t197 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X154 VSS.t125 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X155 VSS VSS.t8 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X156 VSS.t156 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X157 VSS.t218 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X158 VSS.t130 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X159 VSS.t188 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X160 VSS.t145 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X161 VSS VSS.t70 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X162 VSS VSS.t42 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X163 VSS.t216 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X164 VSS.t165 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X165 VSS.t142 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X166 VSS.t121 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X167 VSS.t209 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X168 sky130_asc_nfet_01v8_lvt_1_1/DRAIN vb.t0 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X169 VSS.t170 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X170 VSS.t202 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X171 VSS.t187 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X172 VSS.t169 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X173 sky130_asc_cap_mim_m3_1_4/Cout va.t6 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X174 VSS.t162 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X175 VSS.t207 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X176 VSS.t158 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X177 VDD.t23 VDD.t21 va VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X178 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE.t12 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X179 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_pfet_01v8_lvt_6_1/GATE.t14 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X180 VSS VSS.t22 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X181 VSS.t126 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X182 sky130_asc_nfet_01v8_lvt_1_1/DRAIN va.t0 sky130_asc_cap_mim_m3_1_4/Cout VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X183 va VDD.t18 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X184 VDD.t8 VDD.t6 va VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X185 sky130_asc_pfet_01v8_lvt_6_1/GATE.t7 sky130_asc_pfet_01v8_lvt_6_1/GATE.t6 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X186 VSS.t200 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X187 VSS VSS.t50 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5 area=0p
X188 VSS.t131 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X189 sky130_asc_pfet_01v8_lvt_6_1/GATE vb.t4 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X190 VSS.t160 va sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
R0 VSS.n1631 VSS.n1599 3048.36
R1 VSS.n3836 VSS.n3835 3048.36
R2 VSS.n17829 VSS.n17828 3048.36
R3 VSS.n1139 VSS.n1105 2962.09
R4 VSS.n5102 VSS.n3109 2962.09
R5 VSS.n17902 VSS.n17779 2962.09
R6 VSS.n17854 VSS.n17853 2875.82
R7 VSS.n17878 VSS.n17877 2760.78
R8 VSS.n5137 VSS.n1585 2674.51
R9 VSS.n3811 VSS.n3810 2674.51
R10 VSS.n1163 VSS.n1162 2588.24
R11 VSS.n1162 VSS.n1161 2588.24
R12 VSS.n1161 VSS.n1097 2588.24
R13 VSS.n1155 VSS.n1097 2588.24
R14 VSS.n1155 VSS.n1154 2588.24
R15 VSS.n1154 VSS.n1153 2588.24
R16 VSS.n1153 VSS.n1101 2588.24
R17 VSS.n1147 VSS.n1101 2588.24
R18 VSS.n1147 VSS.n1146 2588.24
R19 VSS.n1146 VSS.n1145 2588.24
R20 VSS.n1145 VSS.n1105 2588.24
R21 VSS.n1121 VSS.n1117 2588.24
R22 VSS.n1122 VSS.n1121 2588.24
R23 VSS.n1123 VSS.n1122 2588.24
R24 VSS.n1123 VSS.n1113 2588.24
R25 VSS.n1129 VSS.n1113 2588.24
R26 VSS.n1130 VSS.n1129 2588.24
R27 VSS.n1131 VSS.n1130 2588.24
R28 VSS.n1131 VSS.n1109 2588.24
R29 VSS.n1137 VSS.n1109 2588.24
R30 VSS.n1138 VSS.n1137 2588.24
R31 VSS.n1139 VSS.n1138 2588.24
R32 VSS.n1318 VSS.n619 2588.24
R33 VSS.n1318 VSS.n1317 2588.24
R34 VSS.n1317 VSS.n1316 2588.24
R35 VSS.n1316 VSS.n626 2588.24
R36 VSS.n1310 VSS.n626 2588.24
R37 VSS.n1310 VSS.n1309 2588.24
R38 VSS.n1309 VSS.n1308 2588.24
R39 VSS.n1308 VSS.n631 2588.24
R40 VSS.n1302 VSS.n631 2588.24
R41 VSS.n1302 VSS.n1301 2588.24
R42 VSS.n1301 VSS.n1300 2588.24
R43 VSS.n1350 VSS.n607 2588.24
R44 VSS.n1344 VSS.n607 2588.24
R45 VSS.n1344 VSS.n1343 2588.24
R46 VSS.n1343 VSS.n1342 2588.24
R47 VSS.n1342 VSS.n611 2588.24
R48 VSS.n1336 VSS.n611 2588.24
R49 VSS.n1336 VSS.n1335 2588.24
R50 VSS.n1335 VSS.n1334 2588.24
R51 VSS.n1334 VSS.n615 2588.24
R52 VSS.n1328 VSS.n615 2588.24
R53 VSS.n1328 VSS.n1327 2588.24
R54 VSS.n5650 VSS.n5649 2588.24
R55 VSS.n5650 VSS.n1359 2588.24
R56 VSS.n5656 VSS.n1359 2588.24
R57 VSS.n5657 VSS.n5656 2588.24
R58 VSS.n5658 VSS.n5657 2588.24
R59 VSS.n5658 VSS.n1355 2588.24
R60 VSS.n5664 VSS.n1355 2588.24
R61 VSS.n5665 VSS.n5664 2588.24
R62 VSS.n5666 VSS.n5665 2588.24
R63 VSS.n5666 VSS.n1351 2588.24
R64 VSS.n5672 VSS.n1351 2588.24
R65 VSS.n1491 VSS.n1462 2588.24
R66 VSS.n1485 VSS.n1462 2588.24
R67 VSS.n1485 VSS.n1484 2588.24
R68 VSS.n1484 VSS.n1483 2588.24
R69 VSS.n1483 VSS.n1466 2588.24
R70 VSS.n1477 VSS.n1466 2588.24
R71 VSS.n1477 VSS.n1476 2588.24
R72 VSS.n1476 VSS.n1475 2588.24
R73 VSS.n1475 VSS.n1470 2588.24
R74 VSS.n1470 VSS.n1364 2588.24
R75 VSS.n5647 VSS.n1364 2588.24
R76 VSS.n5442 VSS.n5441 2588.24
R77 VSS.n5442 VSS.n1500 2588.24
R78 VSS.n5448 VSS.n1500 2588.24
R79 VSS.n5449 VSS.n5448 2588.24
R80 VSS.n5450 VSS.n5449 2588.24
R81 VSS.n5450 VSS.n1496 2588.24
R82 VSS.n5456 VSS.n1496 2588.24
R83 VSS.n5457 VSS.n5456 2588.24
R84 VSS.n5458 VSS.n5457 2588.24
R85 VSS.n5458 VSS.n1492 2588.24
R86 VSS.n5464 VSS.n1492 2588.24
R87 VSS.n1625 VSS.n1599 2588.24
R88 VSS.n1625 VSS.n1624 2588.24
R89 VSS.n1624 VSS.n1623 2588.24
R90 VSS.n1623 VSS.n1603 2588.24
R91 VSS.n1617 VSS.n1603 2588.24
R92 VSS.n1617 VSS.n1616 2588.24
R93 VSS.n1616 VSS.n1615 2588.24
R94 VSS.n1615 VSS.n1607 2588.24
R95 VSS.n1609 VSS.n1607 2588.24
R96 VSS.n1609 VSS.n1505 2588.24
R97 VSS.n5439 VSS.n1505 2588.24
R98 VSS.n1649 VSS.n1588 2588.24
R99 VSS.n1649 VSS.n1648 2588.24
R100 VSS.n1648 VSS.n1647 2588.24
R101 VSS.n1647 VSS.n1590 2588.24
R102 VSS.n1641 VSS.n1590 2588.24
R103 VSS.n1641 VSS.n1640 2588.24
R104 VSS.n1640 VSS.n1639 2588.24
R105 VSS.n1639 VSS.n1595 2588.24
R106 VSS.n1633 VSS.n1595 2588.24
R107 VSS.n1633 VSS.n1632 2588.24
R108 VSS.n1632 VSS.n1631 2588.24
R109 VSS.n5084 VSS.n3121 2588.24
R110 VSS.n5085 VSS.n5084 2588.24
R111 VSS.n5086 VSS.n5085 2588.24
R112 VSS.n5086 VSS.n3117 2588.24
R113 VSS.n5092 VSS.n3117 2588.24
R114 VSS.n5093 VSS.n5092 2588.24
R115 VSS.n5094 VSS.n5093 2588.24
R116 VSS.n5094 VSS.n3113 2588.24
R117 VSS.n5100 VSS.n3113 2588.24
R118 VSS.n5101 VSS.n5100 2588.24
R119 VSS.n5102 VSS.n5101 2588.24
R120 VSS.n5126 VSS.n5125 2588.24
R121 VSS.n5125 VSS.n5124 2588.24
R122 VSS.n5124 VSS.n3101 2588.24
R123 VSS.n5118 VSS.n3101 2588.24
R124 VSS.n5118 VSS.n5117 2588.24
R125 VSS.n5117 VSS.n5116 2588.24
R126 VSS.n5116 VSS.n3105 2588.24
R127 VSS.n5110 VSS.n3105 2588.24
R128 VSS.n5110 VSS.n5109 2588.24
R129 VSS.n5109 VSS.n5108 2588.24
R130 VSS.n5108 VSS.n3109 2588.24
R131 VSS.n5051 VSS.n3136 2588.24
R132 VSS.n5057 VSS.n3136 2588.24
R133 VSS.n5058 VSS.n5057 2588.24
R134 VSS.n5059 VSS.n5058 2588.24
R135 VSS.n5059 VSS.n3132 2588.24
R136 VSS.n5065 VSS.n3132 2588.24
R137 VSS.n5066 VSS.n5065 2588.24
R138 VSS.n5068 VSS.n5066 2588.24
R139 VSS.n5068 VSS.n5067 2588.24
R140 VSS.n5067 VSS.n3128 2588.24
R141 VSS.n5075 VSS.n3128 2588.24
R142 VSS.n3277 VSS.n3243 2588.24
R143 VSS.n3271 VSS.n3243 2588.24
R144 VSS.n3271 VSS.n3270 2588.24
R145 VSS.n3270 VSS.n3269 2588.24
R146 VSS.n3269 VSS.n3247 2588.24
R147 VSS.n3263 VSS.n3247 2588.24
R148 VSS.n3263 VSS.n3262 2588.24
R149 VSS.n3262 VSS.n3261 2588.24
R150 VSS.n3261 VSS.n3251 2588.24
R151 VSS.n3255 VSS.n3251 2588.24
R152 VSS.n3255 VSS.n3140 2588.24
R153 VSS.n4480 VSS.n4479 2588.24
R154 VSS.n4480 VSS.n3286 2588.24
R155 VSS.n4486 VSS.n3286 2588.24
R156 VSS.n4487 VSS.n4486 2588.24
R157 VSS.n4488 VSS.n4487 2588.24
R158 VSS.n4488 VSS.n3282 2588.24
R159 VSS.n4494 VSS.n3282 2588.24
R160 VSS.n4495 VSS.n4494 2588.24
R161 VSS.n4496 VSS.n4495 2588.24
R162 VSS.n4496 VSS.n3278 2588.24
R163 VSS.n4502 VSS.n3278 2588.24
R164 VSS.n4452 VSS.n4451 2588.24
R165 VSS.n4453 VSS.n4452 2588.24
R166 VSS.n4453 VSS.n3301 2588.24
R167 VSS.n4459 VSS.n3301 2588.24
R168 VSS.n4460 VSS.n4459 2588.24
R169 VSS.n4461 VSS.n4460 2588.24
R170 VSS.n4461 VSS.n3297 2588.24
R171 VSS.n4468 VSS.n3297 2588.24
R172 VSS.n4469 VSS.n4468 2588.24
R173 VSS.n4470 VSS.n4469 2588.24
R174 VSS.n4470 VSS.n3290 2588.24
R175 VSS.n3920 VSS.n3887 2588.24
R176 VSS.n3891 VSS.n3887 2588.24
R177 VSS.n3913 VSS.n3891 2588.24
R178 VSS.n3913 VSS.n3912 2588.24
R179 VSS.n3912 VSS.n3911 2588.24
R180 VSS.n3911 VSS.n3892 2588.24
R181 VSS.n3905 VSS.n3892 2588.24
R182 VSS.n3905 VSS.n3904 2588.24
R183 VSS.n3904 VSS.n3903 2588.24
R184 VSS.n3903 VSS.n3896 2588.24
R185 VSS.n3897 VSS.n3896 2588.24
R186 VSS.n3869 VSS.n3417 2588.24
R187 VSS.n3870 VSS.n3869 2588.24
R188 VSS.n3871 VSS.n3870 2588.24
R189 VSS.n3871 VSS.n3413 2588.24
R190 VSS.n3877 VSS.n3413 2588.24
R191 VSS.n3878 VSS.n3877 2588.24
R192 VSS.n3879 VSS.n3878 2588.24
R193 VSS.n3879 VSS.n3409 2588.24
R194 VSS.n3885 VSS.n3409 2588.24
R195 VSS.n3886 VSS.n3885 2588.24
R196 VSS.n3922 VSS.n3886 2588.24
R197 VSS.n3836 VSS.n3432 2588.24
R198 VSS.n3842 VSS.n3432 2588.24
R199 VSS.n3843 VSS.n3842 2588.24
R200 VSS.n3844 VSS.n3843 2588.24
R201 VSS.n3844 VSS.n3428 2588.24
R202 VSS.n3850 VSS.n3428 2588.24
R203 VSS.n3851 VSS.n3850 2588.24
R204 VSS.n3853 VSS.n3851 2588.24
R205 VSS.n3853 VSS.n3852 2588.24
R206 VSS.n3852 VSS.n3424 2588.24
R207 VSS.n3860 VSS.n3424 2588.24
R208 VSS.n3812 VSS.n3444 2588.24
R209 VSS.n3818 VSS.n3444 2588.24
R210 VSS.n3819 VSS.n3818 2588.24
R211 VSS.n3820 VSS.n3819 2588.24
R212 VSS.n3820 VSS.n3440 2588.24
R213 VSS.n3826 VSS.n3440 2588.24
R214 VSS.n3827 VSS.n3826 2588.24
R215 VSS.n3828 VSS.n3827 2588.24
R216 VSS.n3828 VSS.n3436 2588.24
R217 VSS.n3834 VSS.n3436 2588.24
R218 VSS.n3835 VSS.n3834 2588.24
R219 VSS.n17854 VSS.n17803 2588.24
R220 VSS.n17860 VSS.n17803 2588.24
R221 VSS.n17861 VSS.n17860 2588.24
R222 VSS.n17862 VSS.n17861 2588.24
R223 VSS.n17862 VSS.n17799 2588.24
R224 VSS.n17868 VSS.n17799 2588.24
R225 VSS.n17869 VSS.n17868 2588.24
R226 VSS.n17870 VSS.n17869 2588.24
R227 VSS.n17870 VSS.n17795 2588.24
R228 VSS.n17876 VSS.n17795 2588.24
R229 VSS.n17877 VSS.n17876 2588.24
R230 VSS.n17884 VSS.n17791 2588.24
R231 VSS.n17885 VSS.n17884 2588.24
R232 VSS.n17886 VSS.n17885 2588.24
R233 VSS.n17886 VSS.n17787 2588.24
R234 VSS.n17892 VSS.n17787 2588.24
R235 VSS.n17893 VSS.n17892 2588.24
R236 VSS.n17894 VSS.n17893 2588.24
R237 VSS.n17894 VSS.n17783 2588.24
R238 VSS.n17900 VSS.n17783 2588.24
R239 VSS.n17901 VSS.n17900 2588.24
R240 VSS.n17902 VSS.n17901 2588.24
R241 VSS.n17828 VSS.n17827 2588.24
R242 VSS.n17827 VSS.n17822 2588.24
R243 VSS.n17822 VSS.n17774 2588.24
R244 VSS.n17918 VSS.n17774 2588.24
R245 VSS.n17918 VSS.n17917 2588.24
R246 VSS.n17917 VSS.n17916 2588.24
R247 VSS.n17916 VSS.n17775 2588.24
R248 VSS.n17910 VSS.n17775 2588.24
R249 VSS.n17910 VSS.n17909 2588.24
R250 VSS.n17909 VSS.n17908 2588.24
R251 VSS.n17908 VSS.n17779 2588.24
R252 VSS.n17852 VSS.n17808 2588.24
R253 VSS.n17813 VSS.n17808 2588.24
R254 VSS.n17845 VSS.n17813 2588.24
R255 VSS.n17845 VSS.n17844 2588.24
R256 VSS.n17844 VSS.n17843 2588.24
R257 VSS.n17843 VSS.n17814 2588.24
R258 VSS.n17837 VSS.n17814 2588.24
R259 VSS.n17837 VSS.n17836 2588.24
R260 VSS.n17836 VSS.n17835 2588.24
R261 VSS.n17835 VSS.n17818 2588.24
R262 VSS.n17829 VSS.n17818 2588.24
R263 VSS.n1174 VSS.n1092 2473.2
R264 VSS.n4841 VSS.n3100 2473.2
R265 VSS.n1257 VSS.n1256 2099.35
R266 VSS.n1245 VSS.n1026 2099.35
R267 VSS.n1243 VSS.n1035 2099.35
R268 VSS.n1234 VSS.n1233 2099.35
R269 VSS.n1222 VSS.n1045 2099.35
R270 VSS.n1220 VSS.n1054 2099.35
R271 VSS.n1211 VSS.n1210 2099.35
R272 VSS.n1199 VSS.n1064 2099.35
R273 VSS.n1197 VSS.n1073 2099.35
R274 VSS.n1188 VSS.n1187 2099.35
R275 VSS.n1176 VSS.n1083 2099.35
R276 VSS.n929 VSS.n709 2099.35
R277 VSS.n931 VSS.n702 2099.35
R278 VSS.n943 VSS.n942 2099.35
R279 VSS.n953 VSS.n952 2099.35
R280 VSS.n964 VSS.n688 2099.35
R281 VSS.n966 VSS.n681 2099.35
R282 VSS.n978 VSS.n977 2099.35
R283 VSS.n988 VSS.n987 2099.35
R284 VSS.n999 VSS.n667 2099.35
R285 VSS.n1001 VSS.n660 2099.35
R286 VSS.n1013 VSS.n1012 2099.35
R287 VSS.n784 VSS.n774 2099.35
R288 VSS.n796 VSS.n795 2099.35
R289 VSS.n806 VSS.n805 2099.35
R290 VSS.n817 VSS.n760 2099.35
R291 VSS.n819 VSS.n753 2099.35
R292 VSS.n831 VSS.n830 2099.35
R293 VSS.n841 VSS.n840 2099.35
R294 VSS.n852 VSS.n739 2099.35
R295 VSS.n854 VSS.n732 2099.35
R296 VSS.n866 VSS.n865 2099.35
R297 VSS.n876 VSS.n875 2099.35
R298 VSS.n5597 VSS.n5596 2099.35
R299 VSS.n5780 VSS.n5779 2099.35
R300 VSS.n5768 VSS.n526 2099.35
R301 VSS.n5766 VSS.n535 2099.35
R302 VSS.n5757 VSS.n5756 2099.35
R303 VSS.n5745 VSS.n545 2099.35
R304 VSS.n5743 VSS.n554 2099.35
R305 VSS.n5734 VSS.n5733 2099.35
R306 VSS.n5722 VSS.n564 2099.35
R307 VSS.n5720 VSS.n573 2099.35
R308 VSS.n5711 VSS.n5710 2099.35
R309 VSS.n5498 VSS.n1437 2099.35
R310 VSS.n5510 VSS.n5509 2099.35
R311 VSS.n5520 VSS.n5519 2099.35
R312 VSS.n5531 VSS.n1423 2099.35
R313 VSS.n5533 VSS.n1416 2099.35
R314 VSS.n5545 VSS.n5544 2099.35
R315 VSS.n5555 VSS.n5554 2099.35
R316 VSS.n5566 VSS.n1402 2099.35
R317 VSS.n5568 VSS.n1395 2099.35
R318 VSS.n5581 VSS.n5579 2099.35
R319 VSS.n5592 VSS.n1387 2099.35
R320 VSS.n5389 VSS.n5241 2099.35
R321 VSS.n5387 VSS.n5242 2099.35
R322 VSS.n5378 VSS.n5377 2099.35
R323 VSS.n5366 VSS.n5252 2099.35
R324 VSS.n5364 VSS.n5261 2099.35
R325 VSS.n5355 VSS.n5354 2099.35
R326 VSS.n5343 VSS.n5271 2099.35
R327 VSS.n5341 VSS.n5280 2099.35
R328 VSS.n5332 VSS.n5331 2099.35
R329 VSS.n5320 VSS.n5290 2099.35
R330 VSS.n5318 VSS.n5299 2099.35
R331 VSS.n5139 VSS.n1578 2099.35
R332 VSS.n5151 VSS.n5150 2099.35
R333 VSS.n5161 VSS.n5160 2099.35
R334 VSS.n5172 VSS.n1564 2099.35
R335 VSS.n5174 VSS.n1557 2099.35
R336 VSS.n5186 VSS.n5185 2099.35
R337 VSS.n5196 VSS.n5195 2099.35
R338 VSS.n5207 VSS.n1543 2099.35
R339 VSS.n5209 VSS.n1536 2099.35
R340 VSS.n5222 VSS.n5220 2099.35
R341 VSS.n5233 VSS.n1528 2099.35
R342 VSS.n4924 VSS.n4923 2099.35
R343 VSS.n4912 VSS.n4770 2099.35
R344 VSS.n4910 VSS.n4779 2099.35
R345 VSS.n4901 VSS.n4900 2099.35
R346 VSS.n4889 VSS.n4789 2099.35
R347 VSS.n4887 VSS.n4798 2099.35
R348 VSS.n4878 VSS.n4877 2099.35
R349 VSS.n4866 VSS.n4808 2099.35
R350 VSS.n4864 VSS.n4817 2099.35
R351 VSS.n4855 VSS.n4854 2099.35
R352 VSS.n4843 VSS.n4827 2099.35
R353 VSS.n5017 VSS.n5016 2099.35
R354 VSS.n5005 VSS.n4658 2099.35
R355 VSS.n5003 VSS.n4667 2099.35
R356 VSS.n4994 VSS.n4993 2099.35
R357 VSS.n4982 VSS.n4677 2099.35
R358 VSS.n4980 VSS.n4686 2099.35
R359 VSS.n4971 VSS.n4970 2099.35
R360 VSS.n4959 VSS.n4696 2099.35
R361 VSS.n4957 VSS.n4705 2099.35
R362 VSS.n4948 VSS.n4947 2099.35
R363 VSS.n4936 VSS.n4715 2099.35
R364 VSS.n4551 VSS.n4550 2099.35
R365 VSS.n4561 VSS.n4560 2099.35
R366 VSS.n4572 VSS.n3202 2099.35
R367 VSS.n4574 VSS.n3195 2099.35
R368 VSS.n4586 VSS.n4585 2099.35
R369 VSS.n4596 VSS.n4595 2099.35
R370 VSS.n4607 VSS.n3181 2099.35
R371 VSS.n4609 VSS.n3174 2099.35
R372 VSS.n4621 VSS.n4620 2099.35
R373 VSS.n4631 VSS.n4630 2099.35
R374 VSS.n4642 VSS.n3160 2099.35
R375 VSS.n4315 VSS.n4314 2099.35
R376 VSS.n4303 VSS.n4180 2099.35
R377 VSS.n4301 VSS.n4189 2099.35
R378 VSS.n4292 VSS.n4291 2099.35
R379 VSS.n4280 VSS.n4199 2099.35
R380 VSS.n4278 VSS.n4208 2099.35
R381 VSS.n4269 VSS.n4268 2099.35
R382 VSS.n4257 VSS.n4218 2099.35
R383 VSS.n4255 VSS.n4227 2099.35
R384 VSS.n4246 VSS.n4245 2099.35
R385 VSS.n4534 VSS.n3227 2099.35
R386 VSS.n4408 VSS.n4407 2099.35
R387 VSS.n4396 VSS.n4068 2099.35
R388 VSS.n4394 VSS.n4077 2099.35
R389 VSS.n4385 VSS.n4384 2099.35
R390 VSS.n4373 VSS.n4087 2099.35
R391 VSS.n4371 VSS.n4096 2099.35
R392 VSS.n4362 VSS.n4361 2099.35
R393 VSS.n4350 VSS.n4106 2099.35
R394 VSS.n4348 VSS.n4115 2099.35
R395 VSS.n4339 VSS.n4338 2099.35
R396 VSS.n4327 VSS.n4125 2099.35
R397 VSS.n3971 VSS.n3379 2099.35
R398 VSS.n3973 VSS.n3372 2099.35
R399 VSS.n3985 VSS.n3984 2099.35
R400 VSS.n3995 VSS.n3994 2099.35
R401 VSS.n4006 VSS.n3358 2099.35
R402 VSS.n4008 VSS.n3351 2099.35
R403 VSS.n4020 VSS.n4019 2099.35
R404 VSS.n4030 VSS.n4029 2099.35
R405 VSS.n4041 VSS.n3337 2099.35
R406 VSS.n4043 VSS.n3330 2099.35
R407 VSS.n4055 VSS.n4054 2099.35
R408 VSS.n3711 VSS.n3710 2099.35
R409 VSS.n3699 VSS.n3568 2099.35
R410 VSS.n3697 VSS.n3577 2099.35
R411 VSS.n3688 VSS.n3687 2099.35
R412 VSS.n3676 VSS.n3587 2099.35
R413 VSS.n3674 VSS.n3596 2099.35
R414 VSS.n3665 VSS.n3664 2099.35
R415 VSS.n3653 VSS.n3606 2099.35
R416 VSS.n3651 VSS.n3615 2099.35
R417 VSS.n3642 VSS.n3641 2099.35
R418 VSS.n3628 VSS.n3625 2099.35
R419 VSS.n3804 VSS.n3803 2099.35
R420 VSS.n3792 VSS.n3455 2099.35
R421 VSS.n3790 VSS.n3465 2099.35
R422 VSS.n3781 VSS.n3780 2099.35
R423 VSS.n3769 VSS.n3475 2099.35
R424 VSS.n3767 VSS.n3484 2099.35
R425 VSS.n3758 VSS.n3757 2099.35
R426 VSS.n3746 VSS.n3494 2099.35
R427 VSS.n3744 VSS.n3503 2099.35
R428 VSS.n3735 VSS.n3734 2099.35
R429 VSS.n3723 VSS.n3513 2099.35
R430 VSS.n1270 VSS.n648 1294.12
R431 VSS.n1276 VSS.n648 1294.12
R432 VSS.n1277 VSS.n1276 1294.12
R433 VSS.n1278 VSS.n1277 1294.12
R434 VSS.n1278 VSS.n644 1294.12
R435 VSS.n1284 VSS.n644 1294.12
R436 VSS.n1285 VSS.n1284 1294.12
R437 VSS.n1286 VSS.n1285 1294.12
R438 VSS.n1286 VSS.n640 1294.12
R439 VSS.n1292 VSS.n640 1294.12
R440 VSS.n1293 VSS.n1292 1294.12
R441 VSS.n1294 VSS.n1293 1294.12
R442 VSS.n916 VSS.n716 1294.12
R443 VSS.n910 VSS.n716 1294.12
R444 VSS.n910 VSS.n909 1294.12
R445 VSS.n909 VSS.n908 1294.12
R446 VSS.n908 VSS.n888 1294.12
R447 VSS.n902 VSS.n888 1294.12
R448 VSS.n902 VSS.n901 1294.12
R449 VSS.n901 VSS.n900 1294.12
R450 VSS.n900 VSS.n892 1294.12
R451 VSS.n894 VSS.n892 1294.12
R452 VSS.n894 VSS.n620 1294.12
R453 VSS.n1325 VSS.n620 1294.12
R454 VSS.n5698 VSS.n5697 1294.12
R455 VSS.n5697 VSS.n5696 1294.12
R456 VSS.n5696 VSS.n595 1294.12
R457 VSS.n5690 VSS.n595 1294.12
R458 VSS.n5690 VSS.n5689 1294.12
R459 VSS.n5689 VSS.n5688 1294.12
R460 VSS.n5688 VSS.n599 1294.12
R461 VSS.n5682 VSS.n599 1294.12
R462 VSS.n5682 VSS.n5681 1294.12
R463 VSS.n5681 VSS.n5680 1294.12
R464 VSS.n5680 VSS.n603 1294.12
R465 VSS.n5674 VSS.n603 1294.12
R466 VSS.n5621 VSS.n1378 1294.12
R467 VSS.n5622 VSS.n5621 1294.12
R468 VSS.n5623 VSS.n5622 1294.12
R469 VSS.n5623 VSS.n1374 1294.12
R470 VSS.n5629 VSS.n1374 1294.12
R471 VSS.n5630 VSS.n5629 1294.12
R472 VSS.n5631 VSS.n5630 1294.12
R473 VSS.n5631 VSS.n1370 1294.12
R474 VSS.n5638 VSS.n1370 1294.12
R475 VSS.n5639 VSS.n5638 1294.12
R476 VSS.n5640 VSS.n5639 1294.12
R477 VSS.n5640 VSS.n1363 1294.12
R478 VSS.n5490 VSS.n5489 1294.12
R479 VSS.n5489 VSS.n5488 1294.12
R480 VSS.n5488 VSS.n1450 1294.12
R481 VSS.n5482 VSS.n1450 1294.12
R482 VSS.n5482 VSS.n5481 1294.12
R483 VSS.n5481 VSS.n5480 1294.12
R484 VSS.n5480 VSS.n1454 1294.12
R485 VSS.n5474 VSS.n1454 1294.12
R486 VSS.n5474 VSS.n5473 1294.12
R487 VSS.n5473 VSS.n5472 1294.12
R488 VSS.n5472 VSS.n1458 1294.12
R489 VSS.n5466 VSS.n1458 1294.12
R490 VSS.n5413 VSS.n1519 1294.12
R491 VSS.n5414 VSS.n5413 1294.12
R492 VSS.n5415 VSS.n5414 1294.12
R493 VSS.n5415 VSS.n1515 1294.12
R494 VSS.n5421 VSS.n1515 1294.12
R495 VSS.n5422 VSS.n5421 1294.12
R496 VSS.n5423 VSS.n5422 1294.12
R497 VSS.n5423 VSS.n1511 1294.12
R498 VSS.n5430 VSS.n1511 1294.12
R499 VSS.n5431 VSS.n5430 1294.12
R500 VSS.n5432 VSS.n5431 1294.12
R501 VSS.n5432 VSS.n1504 1294.12
R502 VSS.n4757 VSS.n4756 1294.12
R503 VSS.n4756 VSS.n4755 1294.12
R504 VSS.n4755 VSS.n4729 1294.12
R505 VSS.n4749 VSS.n4729 1294.12
R506 VSS.n4749 VSS.n4748 1294.12
R507 VSS.n4748 VSS.n4747 1294.12
R508 VSS.n4747 VSS.n4733 1294.12
R509 VSS.n4741 VSS.n4733 1294.12
R510 VSS.n4741 VSS.n4740 1294.12
R511 VSS.n4740 VSS.n4739 1294.12
R512 VSS.n4739 VSS.n3127 1294.12
R513 VSS.n5077 VSS.n3127 1294.12
R514 VSS.n5026 VSS.n5025 1294.12
R515 VSS.n5027 VSS.n5026 1294.12
R516 VSS.n5027 VSS.n3149 1294.12
R517 VSS.n5033 VSS.n3149 1294.12
R518 VSS.n5034 VSS.n5033 1294.12
R519 VSS.n5035 VSS.n5034 1294.12
R520 VSS.n5035 VSS.n3145 1294.12
R521 VSS.n5041 VSS.n3145 1294.12
R522 VSS.n5042 VSS.n5041 1294.12
R523 VSS.n5043 VSS.n5042 1294.12
R524 VSS.n5043 VSS.n3141 1294.12
R525 VSS.n5049 VSS.n3141 1294.12
R526 VSS.n4528 VSS.n4527 1294.12
R527 VSS.n4527 VSS.n4526 1294.12
R528 VSS.n4526 VSS.n3230 1294.12
R529 VSS.n4520 VSS.n3230 1294.12
R530 VSS.n4520 VSS.n4519 1294.12
R531 VSS.n4519 VSS.n4518 1294.12
R532 VSS.n4518 VSS.n3235 1294.12
R533 VSS.n4512 VSS.n3235 1294.12
R534 VSS.n4512 VSS.n4511 1294.12
R535 VSS.n4511 VSS.n4510 1294.12
R536 VSS.n4510 VSS.n3239 1294.12
R537 VSS.n4504 VSS.n3239 1294.12
R538 VSS.n4167 VSS.n4166 1294.12
R539 VSS.n4166 VSS.n4165 1294.12
R540 VSS.n4165 VSS.n4139 1294.12
R541 VSS.n4159 VSS.n4139 1294.12
R542 VSS.n4159 VSS.n4158 1294.12
R543 VSS.n4158 VSS.n4157 1294.12
R544 VSS.n4157 VSS.n4143 1294.12
R545 VSS.n4151 VSS.n4143 1294.12
R546 VSS.n4151 VSS.n4150 1294.12
R547 VSS.n4150 VSS.n4149 1294.12
R548 VSS.n4149 VSS.n3291 1294.12
R549 VSS.n4477 VSS.n3291 1294.12
R550 VSS.n4421 VSS.n3318 1294.12
R551 VSS.n4427 VSS.n3318 1294.12
R552 VSS.n4428 VSS.n4427 1294.12
R553 VSS.n4429 VSS.n4428 1294.12
R554 VSS.n4429 VSS.n3314 1294.12
R555 VSS.n4435 VSS.n3314 1294.12
R556 VSS.n4436 VSS.n4435 1294.12
R557 VSS.n4437 VSS.n4436 1294.12
R558 VSS.n4437 VSS.n3310 1294.12
R559 VSS.n4443 VSS.n3310 1294.12
R560 VSS.n4444 VSS.n4443 1294.12
R561 VSS.n4445 VSS.n4444 1294.12
R562 VSS.n3947 VSS.n3385 1294.12
R563 VSS.n3947 VSS.n3946 1294.12
R564 VSS.n3946 VSS.n3945 1294.12
R565 VSS.n3945 VSS.n3394 1294.12
R566 VSS.n3939 VSS.n3394 1294.12
R567 VSS.n3939 VSS.n3938 1294.12
R568 VSS.n3938 VSS.n3937 1294.12
R569 VSS.n3937 VSS.n3399 1294.12
R570 VSS.n3931 VSS.n3399 1294.12
R571 VSS.n3931 VSS.n3930 1294.12
R572 VSS.n3930 VSS.n3929 1294.12
R573 VSS.n3929 VSS.n3403 1294.12
R574 VSS.n3555 VSS.n3554 1294.12
R575 VSS.n3554 VSS.n3553 1294.12
R576 VSS.n3553 VSS.n3527 1294.12
R577 VSS.n3547 VSS.n3527 1294.12
R578 VSS.n3547 VSS.n3546 1294.12
R579 VSS.n3546 VSS.n3545 1294.12
R580 VSS.n3545 VSS.n3531 1294.12
R581 VSS.n3539 VSS.n3531 1294.12
R582 VSS.n3539 VSS.n3538 1294.12
R583 VSS.n3538 VSS.n3537 1294.12
R584 VSS.n3537 VSS.n3423 1294.12
R585 VSS.n3862 VSS.n3423 1294.12
R586 VSS.n1294 VSS.n635 1193.46
R587 VSS.n1326 VSS.n1325 1193.46
R588 VSS.n5674 VSS.n5673 1193.46
R589 VSS.n5648 VSS.n1363 1193.46
R590 VSS.n5466 VSS.n5465 1193.46
R591 VSS.n5440 VSS.n1504 1193.46
R592 VSS.n5077 VSS.n5076 1193.46
R593 VSS.n5050 VSS.n5049 1193.46
R594 VSS.n4504 VSS.n4503 1193.46
R595 VSS.n4478 VSS.n4477 1193.46
R596 VSS.n4445 VSS.n3305 1193.46
R597 VSS.n3921 VSS.n3403 1193.46
R598 VSS.n3862 VSS.n3861 1193.46
R599 VSS.n1163 VSS.n1092 1121.57
R600 VSS.n5126 VSS.n3100 1121.57
R601 VSS.n17878 VSS.n17791 1121.57
R602 VSS.n1588 VSS.n1585 1092.81
R603 VSS.n3812 VSS.n3811 1092.81
R604 VSS.n17853 VSS.n17852 1092.81
R605 VSS.n18167 VSS 703.501
R606 VSS.n1117 VSS.n635 690.196
R607 VSS.n1326 VSS.n619 690.196
R608 VSS.n5673 VSS.n1350 690.196
R609 VSS.n5649 VSS.n5648 690.196
R610 VSS.n5465 VSS.n1491 690.196
R611 VSS.n5441 VSS.n5440 690.196
R612 VSS.n5076 VSS.n3121 690.196
R613 VSS.n5051 VSS.n5050 690.196
R614 VSS.n4503 VSS.n3277 690.196
R615 VSS.n4479 VSS.n4478 690.196
R616 VSS.n4451 VSS.n3305 690.196
R617 VSS.n3921 VSS.n3920 690.196
R618 VSS.n3861 VSS.n3417 690.196
R619 VSS.n1178 VSS.n1177 585
R620 VSS.n1177 VSS.n1176 585
R621 VSS.n1085 VSS.n1081 585
R622 VSS.n1187 VSS.n1081 585
R623 VSS.n1077 VSS.n1074 585
R624 VSS.n1074 VSS.n1073 585
R625 VSS.n1201 VSS.n1200 585
R626 VSS.n1200 VSS.n1199 585
R627 VSS.n1066 VSS.n1062 585
R628 VSS.n1210 VSS.n1062 585
R629 VSS.n1058 VSS.n1055 585
R630 VSS.n1055 VSS.n1054 585
R631 VSS.n1224 VSS.n1223 585
R632 VSS.n1223 VSS.n1222 585
R633 VSS.n1047 VSS.n1043 585
R634 VSS.n1233 VSS.n1043 585
R635 VSS.n1039 VSS.n1036 585
R636 VSS.n1036 VSS.n1035 585
R637 VSS.n1247 VSS.n1246 585
R638 VSS.n1246 VSS.n1245 585
R639 VSS.n1028 VSS.n1024 585
R640 VSS.n1256 VSS.n1024 585
R641 VSS.n1022 VSS.n1021 585
R642 VSS.n1022 VSS.n652 585
R643 VSS.n1015 VSS.n1014 585
R644 VSS.n1014 VSS.n1013 585
R645 VSS.n662 VSS.n661 585
R646 VSS.n661 VSS.n660 585
R647 VSS.n998 VSS.n997 585
R648 VSS.n999 VSS.n998 585
R649 VSS.n672 VSS.n671 585
R650 VSS.n988 VSS.n672 585
R651 VSS.n980 VSS.n979 585
R652 VSS.n979 VSS.n978 585
R653 VSS.n683 VSS.n682 585
R654 VSS.n682 VSS.n681 585
R655 VSS.n963 VSS.n962 585
R656 VSS.n964 VSS.n963 585
R657 VSS.n693 VSS.n692 585
R658 VSS.n953 VSS.n693 585
R659 VSS.n945 VSS.n944 585
R660 VSS.n944 VSS.n943 585
R661 VSS.n704 VSS.n703 585
R662 VSS.n703 VSS.n702 585
R663 VSS.n928 VSS.n927 585
R664 VSS.n929 VSS.n928 585
R665 VSS.n714 VSS.n713 585
R666 VSS.n918 VSS.n714 585
R667 VSS.n726 VSS.n722 585
R668 VSS.n876 VSS.n722 585
R669 VSS.n868 VSS.n867 585
R670 VSS.n867 VSS.n866 585
R671 VSS.n734 VSS.n733 585
R672 VSS.n733 VSS.n732 585
R673 VSS.n851 VSS.n850 585
R674 VSS.n852 VSS.n851 585
R675 VSS.n744 VSS.n743 585
R676 VSS.n841 VSS.n744 585
R677 VSS.n833 VSS.n832 585
R678 VSS.n832 VSS.n831 585
R679 VSS.n755 VSS.n754 585
R680 VSS.n754 VSS.n753 585
R681 VSS.n816 VSS.n815 585
R682 VSS.n817 VSS.n816 585
R683 VSS.n765 VSS.n764 585
R684 VSS.n806 VSS.n765 585
R685 VSS.n798 VSS.n797 585
R686 VSS.n797 VSS.n796 585
R687 VSS.n776 VSS.n775 585
R688 VSS.n775 VSS.n774 585
R689 VSS.n781 VSS.n590 585
R690 VSS.n782 VSS.n781 585
R691 VSS.n585 VSS.n581 585
R692 VSS.n5710 VSS.n581 585
R693 VSS.n577 VSS.n574 585
R694 VSS.n574 VSS.n573 585
R695 VSS.n5724 VSS.n5723 585
R696 VSS.n5723 VSS.n5722 585
R697 VSS.n566 VSS.n562 585
R698 VSS.n5733 VSS.n562 585
R699 VSS.n558 VSS.n555 585
R700 VSS.n555 VSS.n554 585
R701 VSS.n5747 VSS.n5746 585
R702 VSS.n5746 VSS.n5745 585
R703 VSS.n547 VSS.n543 585
R704 VSS.n5756 VSS.n543 585
R705 VSS.n539 VSS.n536 585
R706 VSS.n536 VSS.n535 585
R707 VSS.n5770 VSS.n5769 585
R708 VSS.n5769 VSS.n5768 585
R709 VSS.n528 VSS.n524 585
R710 VSS.n5779 VSS.n524 585
R711 VSS.n5599 VSS.n5598 585
R712 VSS.n5598 VSS.n5597 585
R713 VSS.n5607 VSS.n1380 585
R714 VSS.n5608 VSS.n5607 585
R715 VSS.n5591 VSS.n5590 585
R716 VSS.n5592 VSS.n5591 585
R717 VSS.n5583 VSS.n5582 585
R718 VSS.n5582 VSS.n5581 585
R719 VSS.n1397 VSS.n1396 585
R720 VSS.n1396 VSS.n1395 585
R721 VSS.n5565 VSS.n5564 585
R722 VSS.n5566 VSS.n5565 585
R723 VSS.n1407 VSS.n1406 585
R724 VSS.n5555 VSS.n1407 585
R725 VSS.n5547 VSS.n5546 585
R726 VSS.n5546 VSS.n5545 585
R727 VSS.n1418 VSS.n1417 585
R728 VSS.n1417 VSS.n1416 585
R729 VSS.n5530 VSS.n5529 585
R730 VSS.n5531 VSS.n5530 585
R731 VSS.n1428 VSS.n1427 585
R732 VSS.n5520 VSS.n1428 585
R733 VSS.n5512 VSS.n5511 585
R734 VSS.n5511 VSS.n5510 585
R735 VSS.n1439 VSS.n1438 585
R736 VSS.n1438 VSS.n1437 585
R737 VSS.n5495 VSS.n5494 585
R738 VSS.n5496 VSS.n5495 585
R739 VSS.n5304 VSS.n5300 585
R740 VSS.n5300 VSS.n5299 585
R741 VSS.n5322 VSS.n5321 585
R742 VSS.n5321 VSS.n5320 585
R743 VSS.n5292 VSS.n5288 585
R744 VSS.n5331 VSS.n5288 585
R745 VSS.n5284 VSS.n5281 585
R746 VSS.n5281 VSS.n5280 585
R747 VSS.n5345 VSS.n5344 585
R748 VSS.n5344 VSS.n5343 585
R749 VSS.n5273 VSS.n5269 585
R750 VSS.n5354 VSS.n5269 585
R751 VSS.n5265 VSS.n5262 585
R752 VSS.n5262 VSS.n5261 585
R753 VSS.n5368 VSS.n5367 585
R754 VSS.n5367 VSS.n5366 585
R755 VSS.n5254 VSS.n5250 585
R756 VSS.n5377 VSS.n5250 585
R757 VSS.n5246 VSS.n5243 585
R758 VSS.n5243 VSS.n5242 585
R759 VSS.n5391 VSS.n5390 585
R760 VSS.n5390 VSS.n5389 585
R761 VSS.n5399 VSS.n1521 585
R762 VSS.n5400 VSS.n5399 585
R763 VSS.n5232 VSS.n5231 585
R764 VSS.n5233 VSS.n5232 585
R765 VSS.n5224 VSS.n5223 585
R766 VSS.n5223 VSS.n5222 585
R767 VSS.n1538 VSS.n1537 585
R768 VSS.n1537 VSS.n1536 585
R769 VSS.n5206 VSS.n5205 585
R770 VSS.n5207 VSS.n5206 585
R771 VSS.n1548 VSS.n1547 585
R772 VSS.n5196 VSS.n1548 585
R773 VSS.n5188 VSS.n5187 585
R774 VSS.n5187 VSS.n5186 585
R775 VSS.n1559 VSS.n1558 585
R776 VSS.n1558 VSS.n1557 585
R777 VSS.n5171 VSS.n5170 585
R778 VSS.n5172 VSS.n5171 585
R779 VSS.n1569 VSS.n1568 585
R780 VSS.n5161 VSS.n1569 585
R781 VSS.n5153 VSS.n5152 585
R782 VSS.n5152 VSS.n5151 585
R783 VSS.n1580 VSS.n1579 585
R784 VSS.n1579 VSS.n1578 585
R785 VSS.n5136 VSS.n5135 585
R786 VSS.n5137 VSS.n5136 585
R787 VSS.n4845 VSS.n4844 585
R788 VSS.n4844 VSS.n4843 585
R789 VSS.n4829 VSS.n4825 585
R790 VSS.n4854 VSS.n4825 585
R791 VSS.n4821 VSS.n4818 585
R792 VSS.n4818 VSS.n4817 585
R793 VSS.n4868 VSS.n4867 585
R794 VSS.n4867 VSS.n4866 585
R795 VSS.n4810 VSS.n4806 585
R796 VSS.n4877 VSS.n4806 585
R797 VSS.n4802 VSS.n4799 585
R798 VSS.n4799 VSS.n4798 585
R799 VSS.n4891 VSS.n4890 585
R800 VSS.n4890 VSS.n4889 585
R801 VSS.n4791 VSS.n4787 585
R802 VSS.n4900 VSS.n4787 585
R803 VSS.n4783 VSS.n4780 585
R804 VSS.n4780 VSS.n4779 585
R805 VSS.n4914 VSS.n4913 585
R806 VSS.n4913 VSS.n4912 585
R807 VSS.n4772 VSS.n4765 585
R808 VSS.n4923 VSS.n4765 585
R809 VSS.n4767 VSS.n4766 585
R810 VSS.n4768 VSS.n4767 585
R811 VSS.n4938 VSS.n4937 585
R812 VSS.n4937 VSS.n4936 585
R813 VSS.n4717 VSS.n4713 585
R814 VSS.n4947 VSS.n4713 585
R815 VSS.n4709 VSS.n4706 585
R816 VSS.n4706 VSS.n4705 585
R817 VSS.n4961 VSS.n4960 585
R818 VSS.n4960 VSS.n4959 585
R819 VSS.n4698 VSS.n4694 585
R820 VSS.n4970 VSS.n4694 585
R821 VSS.n4690 VSS.n4687 585
R822 VSS.n4687 VSS.n4686 585
R823 VSS.n4984 VSS.n4983 585
R824 VSS.n4983 VSS.n4982 585
R825 VSS.n4679 VSS.n4675 585
R826 VSS.n4993 VSS.n4675 585
R827 VSS.n4671 VSS.n4668 585
R828 VSS.n4668 VSS.n4667 585
R829 VSS.n5007 VSS.n5006 585
R830 VSS.n5006 VSS.n5005 585
R831 VSS.n4660 VSS.n4654 585
R832 VSS.n5016 VSS.n4654 585
R833 VSS.n4655 VSS.n3155 585
R834 VSS.n4656 VSS.n4655 585
R835 VSS.n4641 VSS.n4640 585
R836 VSS.n4642 VSS.n4641 585
R837 VSS.n3165 VSS.n3164 585
R838 VSS.n4631 VSS.n3165 585
R839 VSS.n4623 VSS.n4622 585
R840 VSS.n4622 VSS.n4621 585
R841 VSS.n3176 VSS.n3175 585
R842 VSS.n3175 VSS.n3174 585
R843 VSS.n4606 VSS.n4605 585
R844 VSS.n4607 VSS.n4606 585
R845 VSS.n3186 VSS.n3185 585
R846 VSS.n4596 VSS.n3186 585
R847 VSS.n4588 VSS.n4587 585
R848 VSS.n4587 VSS.n4586 585
R849 VSS.n3197 VSS.n3196 585
R850 VSS.n3196 VSS.n3195 585
R851 VSS.n4571 VSS.n4570 585
R852 VSS.n4572 VSS.n4571 585
R853 VSS.n3207 VSS.n3206 585
R854 VSS.n4561 VSS.n3207 585
R855 VSS.n4553 VSS.n4552 585
R856 VSS.n4552 VSS.n4551 585
R857 VSS.n3218 VSS.n3217 585
R858 VSS.n3217 VSS.n3216 585
R859 VSS.n4536 VSS.n4535 585
R860 VSS.n4535 VSS.n4534 585
R861 VSS.n4237 VSS.n4235 585
R862 VSS.n4245 VSS.n4235 585
R863 VSS.n4231 VSS.n4228 585
R864 VSS.n4228 VSS.n4227 585
R865 VSS.n4259 VSS.n4258 585
R866 VSS.n4258 VSS.n4257 585
R867 VSS.n4220 VSS.n4216 585
R868 VSS.n4268 VSS.n4216 585
R869 VSS.n4212 VSS.n4209 585
R870 VSS.n4209 VSS.n4208 585
R871 VSS.n4282 VSS.n4281 585
R872 VSS.n4281 VSS.n4280 585
R873 VSS.n4201 VSS.n4197 585
R874 VSS.n4291 VSS.n4197 585
R875 VSS.n4193 VSS.n4190 585
R876 VSS.n4190 VSS.n4189 585
R877 VSS.n4305 VSS.n4304 585
R878 VSS.n4304 VSS.n4303 585
R879 VSS.n4182 VSS.n4175 585
R880 VSS.n4314 VSS.n4175 585
R881 VSS.n4177 VSS.n4176 585
R882 VSS.n4178 VSS.n4177 585
R883 VSS.n4329 VSS.n4328 585
R884 VSS.n4328 VSS.n4327 585
R885 VSS.n4127 VSS.n4123 585
R886 VSS.n4338 VSS.n4123 585
R887 VSS.n4119 VSS.n4116 585
R888 VSS.n4116 VSS.n4115 585
R889 VSS.n4352 VSS.n4351 585
R890 VSS.n4351 VSS.n4350 585
R891 VSS.n4108 VSS.n4104 585
R892 VSS.n4361 VSS.n4104 585
R893 VSS.n4100 VSS.n4097 585
R894 VSS.n4097 VSS.n4096 585
R895 VSS.n4375 VSS.n4374 585
R896 VSS.n4374 VSS.n4373 585
R897 VSS.n4089 VSS.n4085 585
R898 VSS.n4384 VSS.n4085 585
R899 VSS.n4081 VSS.n4078 585
R900 VSS.n4078 VSS.n4077 585
R901 VSS.n4398 VSS.n4397 585
R902 VSS.n4397 VSS.n4396 585
R903 VSS.n4070 VSS.n4066 585
R904 VSS.n4407 VSS.n4066 585
R905 VSS.n4064 VSS.n4063 585
R906 VSS.n4064 VSS.n3322 585
R907 VSS.n4057 VSS.n4056 585
R908 VSS.n4056 VSS.n4055 585
R909 VSS.n3332 VSS.n3331 585
R910 VSS.n3331 VSS.n3330 585
R911 VSS.n4040 VSS.n4039 585
R912 VSS.n4041 VSS.n4040 585
R913 VSS.n3342 VSS.n3341 585
R914 VSS.n4030 VSS.n3342 585
R915 VSS.n4022 VSS.n4021 585
R916 VSS.n4021 VSS.n4020 585
R917 VSS.n3353 VSS.n3352 585
R918 VSS.n3352 VSS.n3351 585
R919 VSS.n4005 VSS.n4004 585
R920 VSS.n4006 VSS.n4005 585
R921 VSS.n3363 VSS.n3362 585
R922 VSS.n3995 VSS.n3363 585
R923 VSS.n3987 VSS.n3986 585
R924 VSS.n3986 VSS.n3985 585
R925 VSS.n3374 VSS.n3373 585
R926 VSS.n3373 VSS.n3372 585
R927 VSS.n3970 VSS.n3969 585
R928 VSS.n3971 VSS.n3970 585
R929 VSS.n3384 VSS.n3383 585
R930 VSS.n3960 VSS.n3384 585
R931 VSS.n3630 VSS.n3629 585
R932 VSS.n3629 VSS.n3628 585
R933 VSS.n3627 VSS.n3623 585
R934 VSS.n3641 VSS.n3623 585
R935 VSS.n3619 VSS.n3616 585
R936 VSS.n3616 VSS.n3615 585
R937 VSS.n3655 VSS.n3654 585
R938 VSS.n3654 VSS.n3653 585
R939 VSS.n3608 VSS.n3604 585
R940 VSS.n3664 VSS.n3604 585
R941 VSS.n3600 VSS.n3597 585
R942 VSS.n3597 VSS.n3596 585
R943 VSS.n3678 VSS.n3677 585
R944 VSS.n3677 VSS.n3676 585
R945 VSS.n3589 VSS.n3585 585
R946 VSS.n3687 VSS.n3585 585
R947 VSS.n3581 VSS.n3578 585
R948 VSS.n3578 VSS.n3577 585
R949 VSS.n3701 VSS.n3700 585
R950 VSS.n3700 VSS.n3699 585
R951 VSS.n3570 VSS.n3563 585
R952 VSS.n3710 VSS.n3563 585
R953 VSS.n3565 VSS.n3564 585
R954 VSS.n3566 VSS.n3565 585
R955 VSS.n3725 VSS.n3724 585
R956 VSS.n3724 VSS.n3723 585
R957 VSS.n3515 VSS.n3511 585
R958 VSS.n3734 VSS.n3511 585
R959 VSS.n3507 VSS.n3504 585
R960 VSS.n3504 VSS.n3503 585
R961 VSS.n3748 VSS.n3747 585
R962 VSS.n3747 VSS.n3746 585
R963 VSS.n3496 VSS.n3492 585
R964 VSS.n3757 VSS.n3492 585
R965 VSS.n3488 VSS.n3485 585
R966 VSS.n3485 VSS.n3484 585
R967 VSS.n3771 VSS.n3770 585
R968 VSS.n3770 VSS.n3769 585
R969 VSS.n3477 VSS.n3473 585
R970 VSS.n3780 VSS.n3473 585
R971 VSS.n3469 VSS.n3466 585
R972 VSS.n3466 VSS.n3465 585
R973 VSS.n3794 VSS.n3793 585
R974 VSS.n3793 VSS.n3792 585
R975 VSS.n3457 VSS.n3454 585
R976 VSS.n3803 VSS.n3454 585
R977 VSS.n3809 VSS.n3808 585
R978 VSS.n3810 VSS.n3809 585
R979 VSS.n16336 VSS.n16335 575.163
R980 VSS.n16081 VSS.n16080 575.163
R981 VSS.n15836 VSS.n15835 575.163
R982 VSS.n15593 VSS.n15592 575.163
R983 VSS.n15348 VSS.n15347 575.163
R984 VSS.n15105 VSS.n15104 575.163
R985 VSS.n14860 VSS.n14859 575.163
R986 VSS.n12385 VSS.n12384 575.163
R987 VSS.n12130 VSS.n12129 575.163
R988 VSS.n11885 VSS.n11884 575.163
R989 VSS.n11642 VSS.n11641 575.163
R990 VSS.n11397 VSS.n11396 575.163
R991 VSS.n11154 VSS.n11153 575.163
R992 VSS.n10909 VSS.n10908 575.163
R993 VSS.n8953 VSS.n8952 575.163
R994 VSS.n8698 VSS.n8697 575.163
R995 VSS.n8453 VSS.n8452 575.163
R996 VSS.n8210 VSS.n8209 575.163
R997 VSS.n7965 VSS.n7964 575.163
R998 VSS.n7722 VSS.n7721 575.163
R999 VSS.n7477 VSS.n7476 575.163
R1000 VSS.n1300 VSS.n635 575.163
R1001 VSS.n1327 VSS.n1326 575.163
R1002 VSS.n5673 VSS.n5672 575.163
R1003 VSS.n5648 VSS.n5647 575.163
R1004 VSS.n5465 VSS.n5464 575.163
R1005 VSS.n5440 VSS.n5439 575.163
R1006 VSS.n5076 VSS.n5075 575.163
R1007 VSS.n5050 VSS.n3140 575.163
R1008 VSS.n4503 VSS.n4502 575.163
R1009 VSS.n4478 VSS.n3290 575.163
R1010 VSS.n3897 VSS.n3305 575.163
R1011 VSS.n3922 VSS.n3921 575.163
R1012 VSS.n3861 VSS.n3860 575.163
R1013 VSS.n1269 VSS.n652 488.888
R1014 VSS.n918 VSS.n917 488.888
R1015 VSS.n782 VSS.n594 488.888
R1016 VSS.n5609 VSS.n5608 488.888
R1017 VSS.n5496 VSS.n1444 488.888
R1018 VSS.n5401 VSS.n5400 488.888
R1019 VSS.n4768 VSS.n4724 488.888
R1020 VSS.n4656 VSS.n3153 488.888
R1021 VSS.n3228 VSS.n3216 488.888
R1022 VSS.n4178 VSS.n4134 488.888
R1023 VSS.n4420 VSS.n3322 488.888
R1024 VSS.n3960 VSS.n3959 488.888
R1025 VSS.n3566 VSS.n3522 488.888
R1026 VSS.n1270 VSS.n1269 345.098
R1027 VSS.n917 VSS.n916 345.098
R1028 VSS.n5698 VSS.n594 345.098
R1029 VSS.n5609 VSS.n1378 345.098
R1030 VSS.n5490 VSS.n1444 345.098
R1031 VSS.n5401 VSS.n1519 345.098
R1032 VSS.n4757 VSS.n4724 345.098
R1033 VSS.n5025 VSS.n3153 345.098
R1034 VSS.n4528 VSS.n3228 345.098
R1035 VSS.n4167 VSS.n4134 345.098
R1036 VSS.n4421 VSS.n4420 345.098
R1037 VSS.n3959 VSS.n3385 345.098
R1038 VSS.n3555 VSS.n3522 345.098
R1039 VSS.n14648 VSS.n14647 321.258
R1040 VSS.n10697 VSS.n10696 321.258
R1041 VSS.n7265 VSS.n7264 321.258
R1042 VSS.n1653 VSS.n1585 321.258
R1043 VSS.n3811 VSS.n3448 321.258
R1044 VSS.n17853 VSS.n17807 321.258
R1045 VSS.n14641 VSS.n14640 292.5
R1046 VSS.n14640 VSS.n14639 292.5
R1047 VSS.n14608 VSS.n14607 292.5
R1048 VSS.n14607 VSS.n14606 292.5
R1049 VSS.n14611 VSS.n14610 292.5
R1050 VSS.n14610 VSS.n14609 292.5
R1051 VSS.n14614 VSS.n14613 292.5
R1052 VSS.n14613 VSS.n14612 292.5
R1053 VSS.n14617 VSS.n14616 292.5
R1054 VSS.n14616 VSS.n14615 292.5
R1055 VSS.n14620 VSS.n14619 292.5
R1056 VSS.n14619 VSS.n14618 292.5
R1057 VSS.n14623 VSS.n14622 292.5
R1058 VSS.n14622 VSS.n14621 292.5
R1059 VSS.n14626 VSS.n14625 292.5
R1060 VSS.n14625 VSS.n14624 292.5
R1061 VSS.n14629 VSS.n14628 292.5
R1062 VSS.n14628 VSS.n14627 292.5
R1063 VSS.n14632 VSS.n14631 292.5
R1064 VSS.n14631 VSS.n14630 292.5
R1065 VSS.n14635 VSS.n14634 292.5
R1066 VSS.n14634 VSS.n14633 292.5
R1067 VSS.n14638 VSS.n14637 292.5
R1068 VSS.n14637 VSS.n14636 292.5
R1069 VSS.n16578 VSS.n16577 292.5
R1070 VSS.n16456 VSS.n16455 292.5
R1071 VSS.n16566 VSS.n16565 292.5
R1072 VSS.n16565 VSS.n16564 292.5
R1073 VSS.n16563 VSS.n16562 292.5
R1074 VSS.n16562 VSS.n16561 292.5
R1075 VSS.n16560 VSS.n16559 292.5
R1076 VSS.n16559 VSS.n16558 292.5
R1077 VSS.n16557 VSS.n16556 292.5
R1078 VSS.n16556 VSS.n16555 292.5
R1079 VSS.n16554 VSS.n16553 292.5
R1080 VSS.n16553 VSS.n16552 292.5
R1081 VSS.n16551 VSS.n16550 292.5
R1082 VSS.n16550 VSS.n16549 292.5
R1083 VSS.n16548 VSS.n16547 292.5
R1084 VSS.n16547 VSS.n16546 292.5
R1085 VSS.n16545 VSS.n16544 292.5
R1086 VSS.n16544 VSS.n16543 292.5
R1087 VSS.n16542 VSS.n16541 292.5
R1088 VSS.n16541 VSS.n16540 292.5
R1089 VSS.n16539 VSS.n16538 292.5
R1090 VSS.n16538 VSS.n16537 292.5
R1091 VSS.n16536 VSS.n16535 292.5
R1092 VSS.n16535 VSS.n16534 292.5
R1093 VSS.n16569 VSS.n16568 292.5
R1094 VSS.n16568 VSS.n16567 292.5
R1095 VSS.n16317 VSS.n16316 292.5
R1096 VSS.n16316 VSS.n16315 292.5
R1097 VSS.n16314 VSS.n16313 292.5
R1098 VSS.n16313 VSS.n16312 292.5
R1099 VSS.n16311 VSS.n16310 292.5
R1100 VSS.n16310 VSS.n16309 292.5
R1101 VSS.n16308 VSS.n16307 292.5
R1102 VSS.n16307 VSS.n16306 292.5
R1103 VSS.n16305 VSS.n16304 292.5
R1104 VSS.n16304 VSS.n16303 292.5
R1105 VSS.n16302 VSS.n16301 292.5
R1106 VSS.n16301 VSS.n16300 292.5
R1107 VSS.n16299 VSS.n16298 292.5
R1108 VSS.n16298 VSS.n16297 292.5
R1109 VSS.n16296 VSS.n16295 292.5
R1110 VSS.n16295 VSS.n16294 292.5
R1111 VSS.n16293 VSS.n16292 292.5
R1112 VSS.n16292 VSS.n16291 292.5
R1113 VSS.n16290 VSS.n16289 292.5
R1114 VSS.n16289 VSS.n16288 292.5
R1115 VSS.n16530 VSS.n16529 292.5
R1116 VSS.n16529 VSS.n16528 292.5
R1117 VSS.n16533 VSS.n16532 292.5
R1118 VSS.n16532 VSS.n16531 292.5
R1119 VSS.n16062 VSS.n16061 292.5
R1120 VSS.n16061 VSS.n16060 292.5
R1121 VSS.n16059 VSS.n16058 292.5
R1122 VSS.n16058 VSS.n16057 292.5
R1123 VSS.n16056 VSS.n16055 292.5
R1124 VSS.n16055 VSS.n16054 292.5
R1125 VSS.n16053 VSS.n16052 292.5
R1126 VSS.n16052 VSS.n16051 292.5
R1127 VSS.n16050 VSS.n16049 292.5
R1128 VSS.n16049 VSS.n16048 292.5
R1129 VSS.n16047 VSS.n16046 292.5
R1130 VSS.n16046 VSS.n16045 292.5
R1131 VSS.n16320 VSS.n16319 292.5
R1132 VSS.n16319 VSS.n16318 292.5
R1133 VSS.n16323 VSS.n16322 292.5
R1134 VSS.n16322 VSS.n16321 292.5
R1135 VSS.n16326 VSS.n16325 292.5
R1136 VSS.n16325 VSS.n16324 292.5
R1137 VSS.n16329 VSS.n16328 292.5
R1138 VSS.n16328 VSS.n16327 292.5
R1139 VSS.n16332 VSS.n16331 292.5
R1140 VSS.n16331 VSS.n16330 292.5
R1141 VSS.n16337 VSS.n16336 292.5
R1142 VSS.n16200 VSS.n16199 292.5
R1143 VSS.n15956 VSS.n15955 292.5
R1144 VSS.n15817 VSS.n15816 292.5
R1145 VSS.n15816 VSS.n15815 292.5
R1146 VSS.n15814 VSS.n15813 292.5
R1147 VSS.n15813 VSS.n15812 292.5
R1148 VSS.n15811 VSS.n15810 292.5
R1149 VSS.n15810 VSS.n15809 292.5
R1150 VSS.n15808 VSS.n15807 292.5
R1151 VSS.n15807 VSS.n15806 292.5
R1152 VSS.n15805 VSS.n15804 292.5
R1153 VSS.n15804 VSS.n15803 292.5
R1154 VSS.n15802 VSS.n15801 292.5
R1155 VSS.n15801 VSS.n15800 292.5
R1156 VSS.n16065 VSS.n16064 292.5
R1157 VSS.n16064 VSS.n16063 292.5
R1158 VSS.n16068 VSS.n16067 292.5
R1159 VSS.n16067 VSS.n16066 292.5
R1160 VSS.n16071 VSS.n16070 292.5
R1161 VSS.n16070 VSS.n16069 292.5
R1162 VSS.n16074 VSS.n16073 292.5
R1163 VSS.n16073 VSS.n16072 292.5
R1164 VSS.n16077 VSS.n16076 292.5
R1165 VSS.n16076 VSS.n16075 292.5
R1166 VSS.n16082 VSS.n16081 292.5
R1167 VSS.n15574 VSS.n15573 292.5
R1168 VSS.n15573 VSS.n15572 292.5
R1169 VSS.n15571 VSS.n15570 292.5
R1170 VSS.n15570 VSS.n15569 292.5
R1171 VSS.n15568 VSS.n15567 292.5
R1172 VSS.n15567 VSS.n15566 292.5
R1173 VSS.n15565 VSS.n15564 292.5
R1174 VSS.n15564 VSS.n15563 292.5
R1175 VSS.n15562 VSS.n15561 292.5
R1176 VSS.n15561 VSS.n15560 292.5
R1177 VSS.n15559 VSS.n15558 292.5
R1178 VSS.n15558 VSS.n15557 292.5
R1179 VSS.n15820 VSS.n15819 292.5
R1180 VSS.n15819 VSS.n15818 292.5
R1181 VSS.n15823 VSS.n15822 292.5
R1182 VSS.n15822 VSS.n15821 292.5
R1183 VSS.n15826 VSS.n15825 292.5
R1184 VSS.n15825 VSS.n15824 292.5
R1185 VSS.n15829 VSS.n15828 292.5
R1186 VSS.n15828 VSS.n15827 292.5
R1187 VSS.n15832 VSS.n15831 292.5
R1188 VSS.n15831 VSS.n15830 292.5
R1189 VSS.n15837 VSS.n15836 292.5
R1190 VSS.n15712 VSS.n15711 292.5
R1191 VSS.n15468 VSS.n15467 292.5
R1192 VSS.n15329 VSS.n15328 292.5
R1193 VSS.n15328 VSS.n15327 292.5
R1194 VSS.n15326 VSS.n15325 292.5
R1195 VSS.n15325 VSS.n15324 292.5
R1196 VSS.n15323 VSS.n15322 292.5
R1197 VSS.n15322 VSS.n15321 292.5
R1198 VSS.n15320 VSS.n15319 292.5
R1199 VSS.n15319 VSS.n15318 292.5
R1200 VSS.n15317 VSS.n15316 292.5
R1201 VSS.n15316 VSS.n15315 292.5
R1202 VSS.n15314 VSS.n15313 292.5
R1203 VSS.n15313 VSS.n15312 292.5
R1204 VSS.n15577 VSS.n15576 292.5
R1205 VSS.n15576 VSS.n15575 292.5
R1206 VSS.n15580 VSS.n15579 292.5
R1207 VSS.n15579 VSS.n15578 292.5
R1208 VSS.n15583 VSS.n15582 292.5
R1209 VSS.n15582 VSS.n15581 292.5
R1210 VSS.n15586 VSS.n15585 292.5
R1211 VSS.n15585 VSS.n15584 292.5
R1212 VSS.n15589 VSS.n15588 292.5
R1213 VSS.n15588 VSS.n15587 292.5
R1214 VSS.n15594 VSS.n15593 292.5
R1215 VSS.n15086 VSS.n15085 292.5
R1216 VSS.n15085 VSS.n15084 292.5
R1217 VSS.n15083 VSS.n15082 292.5
R1218 VSS.n15082 VSS.n15081 292.5
R1219 VSS.n15080 VSS.n15079 292.5
R1220 VSS.n15079 VSS.n15078 292.5
R1221 VSS.n15077 VSS.n15076 292.5
R1222 VSS.n15076 VSS.n15075 292.5
R1223 VSS.n15074 VSS.n15073 292.5
R1224 VSS.n15073 VSS.n15072 292.5
R1225 VSS.n15071 VSS.n15070 292.5
R1226 VSS.n15070 VSS.n15069 292.5
R1227 VSS.n15332 VSS.n15331 292.5
R1228 VSS.n15331 VSS.n15330 292.5
R1229 VSS.n15335 VSS.n15334 292.5
R1230 VSS.n15334 VSS.n15333 292.5
R1231 VSS.n15338 VSS.n15337 292.5
R1232 VSS.n15337 VSS.n15336 292.5
R1233 VSS.n15341 VSS.n15340 292.5
R1234 VSS.n15340 VSS.n15339 292.5
R1235 VSS.n15344 VSS.n15343 292.5
R1236 VSS.n15343 VSS.n15342 292.5
R1237 VSS.n15349 VSS.n15348 292.5
R1238 VSS.n15224 VSS.n15223 292.5
R1239 VSS.n14980 VSS.n14979 292.5
R1240 VSS.n14829 VSS.n14828 292.5
R1241 VSS.n14828 VSS.n14827 292.5
R1242 VSS.n14826 VSS.n14825 292.5
R1243 VSS.n14825 VSS.n14824 292.5
R1244 VSS.n14823 VSS.n14822 292.5
R1245 VSS.n14822 VSS.n14821 292.5
R1246 VSS.n14820 VSS.n14819 292.5
R1247 VSS.n14819 VSS.n14818 292.5
R1248 VSS.n14817 VSS.n14816 292.5
R1249 VSS.n14816 VSS.n14815 292.5
R1250 VSS.n14814 VSS.n14813 292.5
R1251 VSS.n14813 VSS.n14812 292.5
R1252 VSS.n15089 VSS.n15088 292.5
R1253 VSS.n15088 VSS.n15087 292.5
R1254 VSS.n15092 VSS.n15091 292.5
R1255 VSS.n15091 VSS.n15090 292.5
R1256 VSS.n15095 VSS.n15094 292.5
R1257 VSS.n15094 VSS.n15093 292.5
R1258 VSS.n15098 VSS.n15097 292.5
R1259 VSS.n15097 VSS.n15096 292.5
R1260 VSS.n15101 VSS.n15100 292.5
R1261 VSS.n15100 VSS.n15099 292.5
R1262 VSS.n15106 VSS.n15105 292.5
R1263 VSS.n14602 VSS.n14601 292.5
R1264 VSS.n14601 VSS.n14600 292.5
R1265 VSS.n14832 VSS.n14831 292.5
R1266 VSS.n14831 VSS.n14830 292.5
R1267 VSS.n14835 VSS.n14834 292.5
R1268 VSS.n14834 VSS.n14833 292.5
R1269 VSS.n14838 VSS.n14837 292.5
R1270 VSS.n14837 VSS.n14836 292.5
R1271 VSS.n14841 VSS.n14840 292.5
R1272 VSS.n14840 VSS.n14839 292.5
R1273 VSS.n14844 VSS.n14843 292.5
R1274 VSS.n14843 VSS.n14842 292.5
R1275 VSS.n14847 VSS.n14846 292.5
R1276 VSS.n14846 VSS.n14845 292.5
R1277 VSS.n14850 VSS.n14849 292.5
R1278 VSS.n14849 VSS.n14848 292.5
R1279 VSS.n14853 VSS.n14852 292.5
R1280 VSS.n14852 VSS.n14851 292.5
R1281 VSS.n14856 VSS.n14855 292.5
R1282 VSS.n14855 VSS.n14854 292.5
R1283 VSS.n14861 VSS.n14860 292.5
R1284 VSS.n14605 VSS.n14604 292.5
R1285 VSS.n14604 VSS.n14603 292.5
R1286 VSS.n14724 VSS.n14723 292.5
R1287 VSS.n10690 VSS.n10689 292.5
R1288 VSS.n10689 VSS.n10688 292.5
R1289 VSS.n10657 VSS.n10656 292.5
R1290 VSS.n10656 VSS.n10655 292.5
R1291 VSS.n10660 VSS.n10659 292.5
R1292 VSS.n10659 VSS.n10658 292.5
R1293 VSS.n10663 VSS.n10662 292.5
R1294 VSS.n10662 VSS.n10661 292.5
R1295 VSS.n10666 VSS.n10665 292.5
R1296 VSS.n10665 VSS.n10664 292.5
R1297 VSS.n10669 VSS.n10668 292.5
R1298 VSS.n10668 VSS.n10667 292.5
R1299 VSS.n10672 VSS.n10671 292.5
R1300 VSS.n10671 VSS.n10670 292.5
R1301 VSS.n10675 VSS.n10674 292.5
R1302 VSS.n10674 VSS.n10673 292.5
R1303 VSS.n10678 VSS.n10677 292.5
R1304 VSS.n10677 VSS.n10676 292.5
R1305 VSS.n10681 VSS.n10680 292.5
R1306 VSS.n10680 VSS.n10679 292.5
R1307 VSS.n10684 VSS.n10683 292.5
R1308 VSS.n10683 VSS.n10682 292.5
R1309 VSS.n10687 VSS.n10686 292.5
R1310 VSS.n10686 VSS.n10685 292.5
R1311 VSS.n12627 VSS.n12626 292.5
R1312 VSS.n12505 VSS.n12504 292.5
R1313 VSS.n12615 VSS.n12614 292.5
R1314 VSS.n12614 VSS.n12613 292.5
R1315 VSS.n12612 VSS.n12611 292.5
R1316 VSS.n12611 VSS.n12610 292.5
R1317 VSS.n12609 VSS.n12608 292.5
R1318 VSS.n12608 VSS.n12607 292.5
R1319 VSS.n12606 VSS.n12605 292.5
R1320 VSS.n12605 VSS.n12604 292.5
R1321 VSS.n12603 VSS.n12602 292.5
R1322 VSS.n12602 VSS.n12601 292.5
R1323 VSS.n12600 VSS.n12599 292.5
R1324 VSS.n12599 VSS.n12598 292.5
R1325 VSS.n12597 VSS.n12596 292.5
R1326 VSS.n12596 VSS.n12595 292.5
R1327 VSS.n12594 VSS.n12593 292.5
R1328 VSS.n12593 VSS.n12592 292.5
R1329 VSS.n12591 VSS.n12590 292.5
R1330 VSS.n12590 VSS.n12589 292.5
R1331 VSS.n12588 VSS.n12587 292.5
R1332 VSS.n12587 VSS.n12586 292.5
R1333 VSS.n12585 VSS.n12584 292.5
R1334 VSS.n12584 VSS.n12583 292.5
R1335 VSS.n12618 VSS.n12617 292.5
R1336 VSS.n12617 VSS.n12616 292.5
R1337 VSS.n12366 VSS.n12365 292.5
R1338 VSS.n12365 VSS.n12364 292.5
R1339 VSS.n12363 VSS.n12362 292.5
R1340 VSS.n12362 VSS.n12361 292.5
R1341 VSS.n12360 VSS.n12359 292.5
R1342 VSS.n12359 VSS.n12358 292.5
R1343 VSS.n12357 VSS.n12356 292.5
R1344 VSS.n12356 VSS.n12355 292.5
R1345 VSS.n12354 VSS.n12353 292.5
R1346 VSS.n12353 VSS.n12352 292.5
R1347 VSS.n12351 VSS.n12350 292.5
R1348 VSS.n12350 VSS.n12349 292.5
R1349 VSS.n12348 VSS.n12347 292.5
R1350 VSS.n12347 VSS.n12346 292.5
R1351 VSS.n12345 VSS.n12344 292.5
R1352 VSS.n12344 VSS.n12343 292.5
R1353 VSS.n12342 VSS.n12341 292.5
R1354 VSS.n12341 VSS.n12340 292.5
R1355 VSS.n12339 VSS.n12338 292.5
R1356 VSS.n12338 VSS.n12337 292.5
R1357 VSS.n12579 VSS.n12578 292.5
R1358 VSS.n12578 VSS.n12577 292.5
R1359 VSS.n12582 VSS.n12581 292.5
R1360 VSS.n12581 VSS.n12580 292.5
R1361 VSS.n12111 VSS.n12110 292.5
R1362 VSS.n12110 VSS.n12109 292.5
R1363 VSS.n12108 VSS.n12107 292.5
R1364 VSS.n12107 VSS.n12106 292.5
R1365 VSS.n12105 VSS.n12104 292.5
R1366 VSS.n12104 VSS.n12103 292.5
R1367 VSS.n12102 VSS.n12101 292.5
R1368 VSS.n12101 VSS.n12100 292.5
R1369 VSS.n12099 VSS.n12098 292.5
R1370 VSS.n12098 VSS.n12097 292.5
R1371 VSS.n12096 VSS.n12095 292.5
R1372 VSS.n12095 VSS.n12094 292.5
R1373 VSS.n12369 VSS.n12368 292.5
R1374 VSS.n12368 VSS.n12367 292.5
R1375 VSS.n12372 VSS.n12371 292.5
R1376 VSS.n12371 VSS.n12370 292.5
R1377 VSS.n12375 VSS.n12374 292.5
R1378 VSS.n12374 VSS.n12373 292.5
R1379 VSS.n12378 VSS.n12377 292.5
R1380 VSS.n12377 VSS.n12376 292.5
R1381 VSS.n12381 VSS.n12380 292.5
R1382 VSS.n12380 VSS.n12379 292.5
R1383 VSS.n12386 VSS.n12385 292.5
R1384 VSS.n12249 VSS.n12248 292.5
R1385 VSS.n12005 VSS.n12004 292.5
R1386 VSS.n11866 VSS.n11865 292.5
R1387 VSS.n11865 VSS.n11864 292.5
R1388 VSS.n11863 VSS.n11862 292.5
R1389 VSS.n11862 VSS.n11861 292.5
R1390 VSS.n11860 VSS.n11859 292.5
R1391 VSS.n11859 VSS.n11858 292.5
R1392 VSS.n11857 VSS.n11856 292.5
R1393 VSS.n11856 VSS.n11855 292.5
R1394 VSS.n11854 VSS.n11853 292.5
R1395 VSS.n11853 VSS.n11852 292.5
R1396 VSS.n11851 VSS.n11850 292.5
R1397 VSS.n11850 VSS.n11849 292.5
R1398 VSS.n12114 VSS.n12113 292.5
R1399 VSS.n12113 VSS.n12112 292.5
R1400 VSS.n12117 VSS.n12116 292.5
R1401 VSS.n12116 VSS.n12115 292.5
R1402 VSS.n12120 VSS.n12119 292.5
R1403 VSS.n12119 VSS.n12118 292.5
R1404 VSS.n12123 VSS.n12122 292.5
R1405 VSS.n12122 VSS.n12121 292.5
R1406 VSS.n12126 VSS.n12125 292.5
R1407 VSS.n12125 VSS.n12124 292.5
R1408 VSS.n12131 VSS.n12130 292.5
R1409 VSS.n11623 VSS.n11622 292.5
R1410 VSS.n11622 VSS.n11621 292.5
R1411 VSS.n11620 VSS.n11619 292.5
R1412 VSS.n11619 VSS.n11618 292.5
R1413 VSS.n11617 VSS.n11616 292.5
R1414 VSS.n11616 VSS.n11615 292.5
R1415 VSS.n11614 VSS.n11613 292.5
R1416 VSS.n11613 VSS.n11612 292.5
R1417 VSS.n11611 VSS.n11610 292.5
R1418 VSS.n11610 VSS.n11609 292.5
R1419 VSS.n11608 VSS.n11607 292.5
R1420 VSS.n11607 VSS.n11606 292.5
R1421 VSS.n11869 VSS.n11868 292.5
R1422 VSS.n11868 VSS.n11867 292.5
R1423 VSS.n11872 VSS.n11871 292.5
R1424 VSS.n11871 VSS.n11870 292.5
R1425 VSS.n11875 VSS.n11874 292.5
R1426 VSS.n11874 VSS.n11873 292.5
R1427 VSS.n11878 VSS.n11877 292.5
R1428 VSS.n11877 VSS.n11876 292.5
R1429 VSS.n11881 VSS.n11880 292.5
R1430 VSS.n11880 VSS.n11879 292.5
R1431 VSS.n11886 VSS.n11885 292.5
R1432 VSS.n11761 VSS.n11760 292.5
R1433 VSS.n11517 VSS.n11516 292.5
R1434 VSS.n11378 VSS.n11377 292.5
R1435 VSS.n11377 VSS.n11376 292.5
R1436 VSS.n11375 VSS.n11374 292.5
R1437 VSS.n11374 VSS.n11373 292.5
R1438 VSS.n11372 VSS.n11371 292.5
R1439 VSS.n11371 VSS.n11370 292.5
R1440 VSS.n11369 VSS.n11368 292.5
R1441 VSS.n11368 VSS.n11367 292.5
R1442 VSS.n11366 VSS.n11365 292.5
R1443 VSS.n11365 VSS.n11364 292.5
R1444 VSS.n11363 VSS.n11362 292.5
R1445 VSS.n11362 VSS.n11361 292.5
R1446 VSS.n11626 VSS.n11625 292.5
R1447 VSS.n11625 VSS.n11624 292.5
R1448 VSS.n11629 VSS.n11628 292.5
R1449 VSS.n11628 VSS.n11627 292.5
R1450 VSS.n11632 VSS.n11631 292.5
R1451 VSS.n11631 VSS.n11630 292.5
R1452 VSS.n11635 VSS.n11634 292.5
R1453 VSS.n11634 VSS.n11633 292.5
R1454 VSS.n11638 VSS.n11637 292.5
R1455 VSS.n11637 VSS.n11636 292.5
R1456 VSS.n11643 VSS.n11642 292.5
R1457 VSS.n11135 VSS.n11134 292.5
R1458 VSS.n11134 VSS.n11133 292.5
R1459 VSS.n11132 VSS.n11131 292.5
R1460 VSS.n11131 VSS.n11130 292.5
R1461 VSS.n11129 VSS.n11128 292.5
R1462 VSS.n11128 VSS.n11127 292.5
R1463 VSS.n11126 VSS.n11125 292.5
R1464 VSS.n11125 VSS.n11124 292.5
R1465 VSS.n11123 VSS.n11122 292.5
R1466 VSS.n11122 VSS.n11121 292.5
R1467 VSS.n11120 VSS.n11119 292.5
R1468 VSS.n11119 VSS.n11118 292.5
R1469 VSS.n11381 VSS.n11380 292.5
R1470 VSS.n11380 VSS.n11379 292.5
R1471 VSS.n11384 VSS.n11383 292.5
R1472 VSS.n11383 VSS.n11382 292.5
R1473 VSS.n11387 VSS.n11386 292.5
R1474 VSS.n11386 VSS.n11385 292.5
R1475 VSS.n11390 VSS.n11389 292.5
R1476 VSS.n11389 VSS.n11388 292.5
R1477 VSS.n11393 VSS.n11392 292.5
R1478 VSS.n11392 VSS.n11391 292.5
R1479 VSS.n11398 VSS.n11397 292.5
R1480 VSS.n11273 VSS.n11272 292.5
R1481 VSS.n11029 VSS.n11028 292.5
R1482 VSS.n10878 VSS.n10877 292.5
R1483 VSS.n10877 VSS.n10876 292.5
R1484 VSS.n10875 VSS.n10874 292.5
R1485 VSS.n10874 VSS.n10873 292.5
R1486 VSS.n10872 VSS.n10871 292.5
R1487 VSS.n10871 VSS.n10870 292.5
R1488 VSS.n10869 VSS.n10868 292.5
R1489 VSS.n10868 VSS.n10867 292.5
R1490 VSS.n10866 VSS.n10865 292.5
R1491 VSS.n10865 VSS.n10864 292.5
R1492 VSS.n10863 VSS.n10862 292.5
R1493 VSS.n10862 VSS.n10861 292.5
R1494 VSS.n11138 VSS.n11137 292.5
R1495 VSS.n11137 VSS.n11136 292.5
R1496 VSS.n11141 VSS.n11140 292.5
R1497 VSS.n11140 VSS.n11139 292.5
R1498 VSS.n11144 VSS.n11143 292.5
R1499 VSS.n11143 VSS.n11142 292.5
R1500 VSS.n11147 VSS.n11146 292.5
R1501 VSS.n11146 VSS.n11145 292.5
R1502 VSS.n11150 VSS.n11149 292.5
R1503 VSS.n11149 VSS.n11148 292.5
R1504 VSS.n11155 VSS.n11154 292.5
R1505 VSS.n10651 VSS.n10650 292.5
R1506 VSS.n10650 VSS.n10649 292.5
R1507 VSS.n10881 VSS.n10880 292.5
R1508 VSS.n10880 VSS.n10879 292.5
R1509 VSS.n10884 VSS.n10883 292.5
R1510 VSS.n10883 VSS.n10882 292.5
R1511 VSS.n10887 VSS.n10886 292.5
R1512 VSS.n10886 VSS.n10885 292.5
R1513 VSS.n10890 VSS.n10889 292.5
R1514 VSS.n10889 VSS.n10888 292.5
R1515 VSS.n10893 VSS.n10892 292.5
R1516 VSS.n10892 VSS.n10891 292.5
R1517 VSS.n10896 VSS.n10895 292.5
R1518 VSS.n10895 VSS.n10894 292.5
R1519 VSS.n10899 VSS.n10898 292.5
R1520 VSS.n10898 VSS.n10897 292.5
R1521 VSS.n10902 VSS.n10901 292.5
R1522 VSS.n10901 VSS.n10900 292.5
R1523 VSS.n10905 VSS.n10904 292.5
R1524 VSS.n10904 VSS.n10903 292.5
R1525 VSS.n10910 VSS.n10909 292.5
R1526 VSS.n10654 VSS.n10653 292.5
R1527 VSS.n10653 VSS.n10652 292.5
R1528 VSS.n10773 VSS.n10772 292.5
R1529 VSS.n7258 VSS.n7257 292.5
R1530 VSS.n7257 VSS.n7256 292.5
R1531 VSS.n7225 VSS.n7224 292.5
R1532 VSS.n7224 VSS.n7223 292.5
R1533 VSS.n7228 VSS.n7227 292.5
R1534 VSS.n7227 VSS.n7226 292.5
R1535 VSS.n7231 VSS.n7230 292.5
R1536 VSS.n7230 VSS.n7229 292.5
R1537 VSS.n7234 VSS.n7233 292.5
R1538 VSS.n7233 VSS.n7232 292.5
R1539 VSS.n7237 VSS.n7236 292.5
R1540 VSS.n7236 VSS.n7235 292.5
R1541 VSS.n7240 VSS.n7239 292.5
R1542 VSS.n7239 VSS.n7238 292.5
R1543 VSS.n7243 VSS.n7242 292.5
R1544 VSS.n7242 VSS.n7241 292.5
R1545 VSS.n7246 VSS.n7245 292.5
R1546 VSS.n7245 VSS.n7244 292.5
R1547 VSS.n7249 VSS.n7248 292.5
R1548 VSS.n7248 VSS.n7247 292.5
R1549 VSS.n7252 VSS.n7251 292.5
R1550 VSS.n7251 VSS.n7250 292.5
R1551 VSS.n7255 VSS.n7254 292.5
R1552 VSS.n7254 VSS.n7253 292.5
R1553 VSS.n9195 VSS.n9194 292.5
R1554 VSS.n9073 VSS.n9072 292.5
R1555 VSS.n9183 VSS.n9182 292.5
R1556 VSS.n9182 VSS.n9181 292.5
R1557 VSS.n9180 VSS.n9179 292.5
R1558 VSS.n9179 VSS.n9178 292.5
R1559 VSS.n9177 VSS.n9176 292.5
R1560 VSS.n9176 VSS.n9175 292.5
R1561 VSS.n9174 VSS.n9173 292.5
R1562 VSS.n9173 VSS.n9172 292.5
R1563 VSS.n9171 VSS.n9170 292.5
R1564 VSS.n9170 VSS.n9169 292.5
R1565 VSS.n9168 VSS.n9167 292.5
R1566 VSS.n9167 VSS.n9166 292.5
R1567 VSS.n9165 VSS.n9164 292.5
R1568 VSS.n9164 VSS.n9163 292.5
R1569 VSS.n9162 VSS.n9161 292.5
R1570 VSS.n9161 VSS.n9160 292.5
R1571 VSS.n9159 VSS.n9158 292.5
R1572 VSS.n9158 VSS.n9157 292.5
R1573 VSS.n9156 VSS.n9155 292.5
R1574 VSS.n9155 VSS.n9154 292.5
R1575 VSS.n9153 VSS.n9152 292.5
R1576 VSS.n9152 VSS.n9151 292.5
R1577 VSS.n9186 VSS.n9185 292.5
R1578 VSS.n9185 VSS.n9184 292.5
R1579 VSS.n8934 VSS.n8933 292.5
R1580 VSS.n8933 VSS.n8932 292.5
R1581 VSS.n8931 VSS.n8930 292.5
R1582 VSS.n8930 VSS.n8929 292.5
R1583 VSS.n8928 VSS.n8927 292.5
R1584 VSS.n8927 VSS.n8926 292.5
R1585 VSS.n8925 VSS.n8924 292.5
R1586 VSS.n8924 VSS.n8923 292.5
R1587 VSS.n8922 VSS.n8921 292.5
R1588 VSS.n8921 VSS.n8920 292.5
R1589 VSS.n8919 VSS.n8918 292.5
R1590 VSS.n8918 VSS.n8917 292.5
R1591 VSS.n8916 VSS.n8915 292.5
R1592 VSS.n8915 VSS.n8914 292.5
R1593 VSS.n8913 VSS.n8912 292.5
R1594 VSS.n8912 VSS.n8911 292.5
R1595 VSS.n8910 VSS.n8909 292.5
R1596 VSS.n8909 VSS.n8908 292.5
R1597 VSS.n8907 VSS.n8906 292.5
R1598 VSS.n8906 VSS.n8905 292.5
R1599 VSS.n9147 VSS.n9146 292.5
R1600 VSS.n9146 VSS.n9145 292.5
R1601 VSS.n9150 VSS.n9149 292.5
R1602 VSS.n9149 VSS.n9148 292.5
R1603 VSS.n8679 VSS.n8678 292.5
R1604 VSS.n8678 VSS.n8677 292.5
R1605 VSS.n8676 VSS.n8675 292.5
R1606 VSS.n8675 VSS.n8674 292.5
R1607 VSS.n8673 VSS.n8672 292.5
R1608 VSS.n8672 VSS.n8671 292.5
R1609 VSS.n8670 VSS.n8669 292.5
R1610 VSS.n8669 VSS.n8668 292.5
R1611 VSS.n8667 VSS.n8666 292.5
R1612 VSS.n8666 VSS.n8665 292.5
R1613 VSS.n8664 VSS.n8663 292.5
R1614 VSS.n8663 VSS.n8662 292.5
R1615 VSS.n8937 VSS.n8936 292.5
R1616 VSS.n8936 VSS.n8935 292.5
R1617 VSS.n8940 VSS.n8939 292.5
R1618 VSS.n8939 VSS.n8938 292.5
R1619 VSS.n8943 VSS.n8942 292.5
R1620 VSS.n8942 VSS.n8941 292.5
R1621 VSS.n8946 VSS.n8945 292.5
R1622 VSS.n8945 VSS.n8944 292.5
R1623 VSS.n8949 VSS.n8948 292.5
R1624 VSS.n8948 VSS.n8947 292.5
R1625 VSS.n8954 VSS.n8953 292.5
R1626 VSS.n8817 VSS.n8816 292.5
R1627 VSS.n8573 VSS.n8572 292.5
R1628 VSS.n8434 VSS.n8433 292.5
R1629 VSS.n8433 VSS.n8432 292.5
R1630 VSS.n8431 VSS.n8430 292.5
R1631 VSS.n8430 VSS.n8429 292.5
R1632 VSS.n8428 VSS.n8427 292.5
R1633 VSS.n8427 VSS.n8426 292.5
R1634 VSS.n8425 VSS.n8424 292.5
R1635 VSS.n8424 VSS.n8423 292.5
R1636 VSS.n8422 VSS.n8421 292.5
R1637 VSS.n8421 VSS.n8420 292.5
R1638 VSS.n8419 VSS.n8418 292.5
R1639 VSS.n8418 VSS.n8417 292.5
R1640 VSS.n8682 VSS.n8681 292.5
R1641 VSS.n8681 VSS.n8680 292.5
R1642 VSS.n8685 VSS.n8684 292.5
R1643 VSS.n8684 VSS.n8683 292.5
R1644 VSS.n8688 VSS.n8687 292.5
R1645 VSS.n8687 VSS.n8686 292.5
R1646 VSS.n8691 VSS.n8690 292.5
R1647 VSS.n8690 VSS.n8689 292.5
R1648 VSS.n8694 VSS.n8693 292.5
R1649 VSS.n8693 VSS.n8692 292.5
R1650 VSS.n8699 VSS.n8698 292.5
R1651 VSS.n8191 VSS.n8190 292.5
R1652 VSS.n8190 VSS.n8189 292.5
R1653 VSS.n8188 VSS.n8187 292.5
R1654 VSS.n8187 VSS.n8186 292.5
R1655 VSS.n8185 VSS.n8184 292.5
R1656 VSS.n8184 VSS.n8183 292.5
R1657 VSS.n8182 VSS.n8181 292.5
R1658 VSS.n8181 VSS.n8180 292.5
R1659 VSS.n8179 VSS.n8178 292.5
R1660 VSS.n8178 VSS.n8177 292.5
R1661 VSS.n8176 VSS.n8175 292.5
R1662 VSS.n8175 VSS.n8174 292.5
R1663 VSS.n8437 VSS.n8436 292.5
R1664 VSS.n8436 VSS.n8435 292.5
R1665 VSS.n8440 VSS.n8439 292.5
R1666 VSS.n8439 VSS.n8438 292.5
R1667 VSS.n8443 VSS.n8442 292.5
R1668 VSS.n8442 VSS.n8441 292.5
R1669 VSS.n8446 VSS.n8445 292.5
R1670 VSS.n8445 VSS.n8444 292.5
R1671 VSS.n8449 VSS.n8448 292.5
R1672 VSS.n8448 VSS.n8447 292.5
R1673 VSS.n8454 VSS.n8453 292.5
R1674 VSS.n8329 VSS.n8328 292.5
R1675 VSS.n8085 VSS.n8084 292.5
R1676 VSS.n7946 VSS.n7945 292.5
R1677 VSS.n7945 VSS.n7944 292.5
R1678 VSS.n7943 VSS.n7942 292.5
R1679 VSS.n7942 VSS.n7941 292.5
R1680 VSS.n7940 VSS.n7939 292.5
R1681 VSS.n7939 VSS.n7938 292.5
R1682 VSS.n7937 VSS.n7936 292.5
R1683 VSS.n7936 VSS.n7935 292.5
R1684 VSS.n7934 VSS.n7933 292.5
R1685 VSS.n7933 VSS.n7932 292.5
R1686 VSS.n7931 VSS.n7930 292.5
R1687 VSS.n7930 VSS.n7929 292.5
R1688 VSS.n8194 VSS.n8193 292.5
R1689 VSS.n8193 VSS.n8192 292.5
R1690 VSS.n8197 VSS.n8196 292.5
R1691 VSS.n8196 VSS.n8195 292.5
R1692 VSS.n8200 VSS.n8199 292.5
R1693 VSS.n8199 VSS.n8198 292.5
R1694 VSS.n8203 VSS.n8202 292.5
R1695 VSS.n8202 VSS.n8201 292.5
R1696 VSS.n8206 VSS.n8205 292.5
R1697 VSS.n8205 VSS.n8204 292.5
R1698 VSS.n8211 VSS.n8210 292.5
R1699 VSS.n7703 VSS.n7702 292.5
R1700 VSS.n7702 VSS.n7701 292.5
R1701 VSS.n7700 VSS.n7699 292.5
R1702 VSS.n7699 VSS.n7698 292.5
R1703 VSS.n7697 VSS.n7696 292.5
R1704 VSS.n7696 VSS.n7695 292.5
R1705 VSS.n7694 VSS.n7693 292.5
R1706 VSS.n7693 VSS.n7692 292.5
R1707 VSS.n7691 VSS.n7690 292.5
R1708 VSS.n7690 VSS.n7689 292.5
R1709 VSS.n7688 VSS.n7687 292.5
R1710 VSS.n7687 VSS.n7686 292.5
R1711 VSS.n7949 VSS.n7948 292.5
R1712 VSS.n7948 VSS.n7947 292.5
R1713 VSS.n7952 VSS.n7951 292.5
R1714 VSS.n7951 VSS.n7950 292.5
R1715 VSS.n7955 VSS.n7954 292.5
R1716 VSS.n7954 VSS.n7953 292.5
R1717 VSS.n7958 VSS.n7957 292.5
R1718 VSS.n7957 VSS.n7956 292.5
R1719 VSS.n7961 VSS.n7960 292.5
R1720 VSS.n7960 VSS.n7959 292.5
R1721 VSS.n7966 VSS.n7965 292.5
R1722 VSS.n7841 VSS.n7840 292.5
R1723 VSS.n7597 VSS.n7596 292.5
R1724 VSS.n7446 VSS.n7445 292.5
R1725 VSS.n7445 VSS.n7444 292.5
R1726 VSS.n7443 VSS.n7442 292.5
R1727 VSS.n7442 VSS.n7441 292.5
R1728 VSS.n7440 VSS.n7439 292.5
R1729 VSS.n7439 VSS.n7438 292.5
R1730 VSS.n7437 VSS.n7436 292.5
R1731 VSS.n7436 VSS.n7435 292.5
R1732 VSS.n7434 VSS.n7433 292.5
R1733 VSS.n7433 VSS.n7432 292.5
R1734 VSS.n7431 VSS.n7430 292.5
R1735 VSS.n7430 VSS.n7429 292.5
R1736 VSS.n7706 VSS.n7705 292.5
R1737 VSS.n7705 VSS.n7704 292.5
R1738 VSS.n7709 VSS.n7708 292.5
R1739 VSS.n7708 VSS.n7707 292.5
R1740 VSS.n7712 VSS.n7711 292.5
R1741 VSS.n7711 VSS.n7710 292.5
R1742 VSS.n7715 VSS.n7714 292.5
R1743 VSS.n7714 VSS.n7713 292.5
R1744 VSS.n7718 VSS.n7717 292.5
R1745 VSS.n7717 VSS.n7716 292.5
R1746 VSS.n7723 VSS.n7722 292.5
R1747 VSS.n7219 VSS.n7218 292.5
R1748 VSS.n7218 VSS.n7217 292.5
R1749 VSS.n7449 VSS.n7448 292.5
R1750 VSS.n7448 VSS.n7447 292.5
R1751 VSS.n7452 VSS.n7451 292.5
R1752 VSS.n7451 VSS.n7450 292.5
R1753 VSS.n7455 VSS.n7454 292.5
R1754 VSS.n7454 VSS.n7453 292.5
R1755 VSS.n7458 VSS.n7457 292.5
R1756 VSS.n7457 VSS.n7456 292.5
R1757 VSS.n7461 VSS.n7460 292.5
R1758 VSS.n7460 VSS.n7459 292.5
R1759 VSS.n7464 VSS.n7463 292.5
R1760 VSS.n7463 VSS.n7462 292.5
R1761 VSS.n7467 VSS.n7466 292.5
R1762 VSS.n7466 VSS.n7465 292.5
R1763 VSS.n7470 VSS.n7469 292.5
R1764 VSS.n7469 VSS.n7468 292.5
R1765 VSS.n7473 VSS.n7472 292.5
R1766 VSS.n7472 VSS.n7471 292.5
R1767 VSS.n7478 VSS.n7477 292.5
R1768 VSS.n7222 VSS.n7221 292.5
R1769 VSS.n7221 VSS.n7220 292.5
R1770 VSS.n7341 VSS.n7340 292.5
R1771 VSS.n1652 VSS.n1651 292.5
R1772 VSS.n1651 VSS.n1588 292.5
R1773 VSS.n1630 VSS.n1629 292.5
R1774 VSS.n1631 VSS.n1630 292.5
R1775 VSS.n1598 VSS.n1597 292.5
R1776 VSS.n1632 VSS.n1598 292.5
R1777 VSS.n1635 VSS.n1634 292.5
R1778 VSS.n1634 VSS.n1633 292.5
R1779 VSS.n1636 VSS.n1596 292.5
R1780 VSS.n1596 VSS.n1595 292.5
R1781 VSS.n1638 VSS.n1637 292.5
R1782 VSS.n1639 VSS.n1638 292.5
R1783 VSS.n1594 VSS.n1593 292.5
R1784 VSS.n1640 VSS.n1594 292.5
R1785 VSS.n1643 VSS.n1642 292.5
R1786 VSS.n1642 VSS.n1641 292.5
R1787 VSS.n1644 VSS.n1591 292.5
R1788 VSS.n1591 VSS.n1590 292.5
R1789 VSS.n1646 VSS.n1645 292.5
R1790 VSS.n1647 VSS.n1646 292.5
R1791 VSS.n1592 VSS.n1589 292.5
R1792 VSS.n1648 VSS.n1589 292.5
R1793 VSS.n1650 VSS.n1587 292.5
R1794 VSS.n1650 VSS.n1649 292.5
R1795 VSS.n1141 VSS.n1140 292.5
R1796 VSS.n1140 VSS.n1139 292.5
R1797 VSS.n1118 VSS.n637 292.5
R1798 VSS.n1118 VSS.n1117 292.5
R1799 VSS.n1120 VSS.n1119 292.5
R1800 VSS.n1121 VSS.n1120 292.5
R1801 VSS.n1116 VSS.n1115 292.5
R1802 VSS.n1122 VSS.n1116 292.5
R1803 VSS.n1125 VSS.n1124 292.5
R1804 VSS.n1124 VSS.n1123 292.5
R1805 VSS.n1126 VSS.n1114 292.5
R1806 VSS.n1114 VSS.n1113 292.5
R1807 VSS.n1128 VSS.n1127 292.5
R1808 VSS.n1129 VSS.n1128 292.5
R1809 VSS.n1112 VSS.n1111 292.5
R1810 VSS.n1130 VSS.n1112 292.5
R1811 VSS.n1133 VSS.n1132 292.5
R1812 VSS.n1132 VSS.n1131 292.5
R1813 VSS.n1134 VSS.n1110 292.5
R1814 VSS.n1110 VSS.n1109 292.5
R1815 VSS.n1136 VSS.n1135 292.5
R1816 VSS.n1137 VSS.n1136 292.5
R1817 VSS.n1108 VSS.n1107 292.5
R1818 VSS.n1138 VSS.n1108 292.5
R1819 VSS.n1096 VSS.n1095 292.5
R1820 VSS.n1162 VSS.n1096 292.5
R1821 VSS.n1160 VSS.n1159 292.5
R1822 VSS.n1161 VSS.n1160 292.5
R1823 VSS.n1158 VSS.n1098 292.5
R1824 VSS.n1098 VSS.n1097 292.5
R1825 VSS.n1157 VSS.n1156 292.5
R1826 VSS.n1156 VSS.n1155 292.5
R1827 VSS.n1100 VSS.n1099 292.5
R1828 VSS.n1154 VSS.n1100 292.5
R1829 VSS.n1152 VSS.n1151 292.5
R1830 VSS.n1153 VSS.n1152 292.5
R1831 VSS.n1150 VSS.n1102 292.5
R1832 VSS.n1102 VSS.n1101 292.5
R1833 VSS.n1149 VSS.n1148 292.5
R1834 VSS.n1148 VSS.n1147 292.5
R1835 VSS.n1104 VSS.n1103 292.5
R1836 VSS.n1146 VSS.n1104 292.5
R1837 VSS.n1144 VSS.n1143 292.5
R1838 VSS.n1145 VSS.n1144 292.5
R1839 VSS.n1142 VSS.n1106 292.5
R1840 VSS.n1106 VSS.n1105 292.5
R1841 VSS.n1165 VSS.n1164 292.5
R1842 VSS.n1164 VSS.n1163 292.5
R1843 VSS.n1166 VSS.n1093 292.5
R1844 VSS.n1093 VSS.n1092 292.5
R1845 VSS.n1023 VSS.n1019 292.5
R1846 VSS.n1025 VSS.n1023 292.5
R1847 VSS.n1254 VSS.n1253 292.5
R1848 VSS.n1255 VSS.n1254 292.5
R1849 VSS.n1034 VSS.n1033 292.5
R1850 VSS.n1244 VSS.n1034 292.5
R1851 VSS.n1042 VSS.n1040 292.5
R1852 VSS.n1044 VSS.n1042 292.5
R1853 VSS.n1231 VSS.n1230 292.5
R1854 VSS.n1232 VSS.n1231 292.5
R1855 VSS.n1053 VSS.n1052 292.5
R1856 VSS.n1221 VSS.n1053 292.5
R1857 VSS.n1061 VSS.n1059 292.5
R1858 VSS.n1063 VSS.n1061 292.5
R1859 VSS.n1208 VSS.n1207 292.5
R1860 VSS.n1209 VSS.n1208 292.5
R1861 VSS.n1072 VSS.n1071 292.5
R1862 VSS.n1198 VSS.n1072 292.5
R1863 VSS.n1080 VSS.n1078 292.5
R1864 VSS.n1082 VSS.n1080 292.5
R1865 VSS.n1185 VSS.n1184 292.5
R1866 VSS.n1186 VSS.n1185 292.5
R1867 VSS.n1091 VSS.n1090 292.5
R1868 VSS.n1175 VSS.n1091 292.5
R1869 VSS.n655 VSS.n654 292.5
R1870 VSS.n654 VSS.n653 292.5
R1871 VSS.n1010 VSS.n1009 292.5
R1872 VSS.n1011 VSS.n1010 292.5
R1873 VSS.n666 VSS.n664 292.5
R1874 VSS.n1000 VSS.n666 292.5
R1875 VSS.n991 VSS.n990 292.5
R1876 VSS.n990 VSS.n989 292.5
R1877 VSS.n675 VSS.n674 292.5
R1878 VSS.n674 VSS.n673 292.5
R1879 VSS.n975 VSS.n974 292.5
R1880 VSS.n976 VSS.n975 292.5
R1881 VSS.n687 VSS.n685 292.5
R1882 VSS.n965 VSS.n687 292.5
R1883 VSS.n956 VSS.n955 292.5
R1884 VSS.n955 VSS.n954 292.5
R1885 VSS.n696 VSS.n695 292.5
R1886 VSS.n695 VSS.n694 292.5
R1887 VSS.n940 VSS.n939 292.5
R1888 VSS.n941 VSS.n940 292.5
R1889 VSS.n708 VSS.n706 292.5
R1890 VSS.n930 VSS.n708 292.5
R1891 VSS.n921 VSS.n920 292.5
R1892 VSS.n920 VSS.n919 292.5
R1893 VSS.n1321 VSS.n1320 292.5
R1894 VSS.n1320 VSS.n619 292.5
R1895 VSS.n1319 VSS.n624 292.5
R1896 VSS.n1319 VSS.n1318 292.5
R1897 VSS.n628 VSS.n625 292.5
R1898 VSS.n1317 VSS.n625 292.5
R1899 VSS.n1315 VSS.n1314 292.5
R1900 VSS.n1316 VSS.n1315 292.5
R1901 VSS.n1313 VSS.n627 292.5
R1902 VSS.n627 VSS.n626 292.5
R1903 VSS.n1312 VSS.n1311 292.5
R1904 VSS.n1311 VSS.n1310 292.5
R1905 VSS.n630 VSS.n629 292.5
R1906 VSS.n1309 VSS.n630 292.5
R1907 VSS.n1307 VSS.n1306 292.5
R1908 VSS.n1308 VSS.n1307 292.5
R1909 VSS.n1305 VSS.n632 292.5
R1910 VSS.n632 VSS.n631 292.5
R1911 VSS.n1304 VSS.n1303 292.5
R1912 VSS.n1303 VSS.n1302 292.5
R1913 VSS.n634 VSS.n633 292.5
R1914 VSS.n1301 VSS.n634 292.5
R1915 VSS.n1299 VSS.n1298 292.5
R1916 VSS.n1300 VSS.n1299 292.5
R1917 VSS.n1349 VSS.n1348 292.5
R1918 VSS.n1350 VSS.n1349 292.5
R1919 VSS.n1347 VSS.n608 292.5
R1920 VSS.n608 VSS.n607 292.5
R1921 VSS.n1346 VSS.n1345 292.5
R1922 VSS.n1345 VSS.n1344 292.5
R1923 VSS.n610 VSS.n609 292.5
R1924 VSS.n1343 VSS.n610 292.5
R1925 VSS.n1341 VSS.n1340 292.5
R1926 VSS.n1342 VSS.n1341 292.5
R1927 VSS.n1339 VSS.n612 292.5
R1928 VSS.n612 VSS.n611 292.5
R1929 VSS.n1338 VSS.n1337 292.5
R1930 VSS.n1337 VSS.n1336 292.5
R1931 VSS.n614 VSS.n613 292.5
R1932 VSS.n1335 VSS.n614 292.5
R1933 VSS.n1333 VSS.n1332 292.5
R1934 VSS.n1334 VSS.n1333 292.5
R1935 VSS.n1331 VSS.n616 292.5
R1936 VSS.n616 VSS.n615 292.5
R1937 VSS.n1330 VSS.n1329 292.5
R1938 VSS.n1329 VSS.n1328 292.5
R1939 VSS.n618 VSS.n617 292.5
R1940 VSS.n1327 VSS.n618 292.5
R1941 VSS.n878 VSS.n721 292.5
R1942 VSS.n878 VSS.n877 292.5
R1943 VSS.n725 VSS.n724 292.5
R1944 VSS.n724 VSS.n723 292.5
R1945 VSS.n863 VSS.n862 292.5
R1946 VSS.n864 VSS.n863 292.5
R1947 VSS.n738 VSS.n736 292.5
R1948 VSS.n853 VSS.n738 292.5
R1949 VSS.n844 VSS.n843 292.5
R1950 VSS.n843 VSS.n842 292.5
R1951 VSS.n747 VSS.n746 292.5
R1952 VSS.n746 VSS.n745 292.5
R1953 VSS.n828 VSS.n827 292.5
R1954 VSS.n829 VSS.n828 292.5
R1955 VSS.n759 VSS.n757 292.5
R1956 VSS.n818 VSS.n759 292.5
R1957 VSS.n809 VSS.n808 292.5
R1958 VSS.n808 VSS.n807 292.5
R1959 VSS.n768 VSS.n767 292.5
R1960 VSS.n767 VSS.n766 292.5
R1961 VSS.n793 VSS.n792 292.5
R1962 VSS.n794 VSS.n793 292.5
R1963 VSS.n780 VSS.n778 292.5
R1964 VSS.n783 VSS.n780 292.5
R1965 VSS.n5708 VSS.n5707 292.5
R1966 VSS.n5709 VSS.n5708 292.5
R1967 VSS.n580 VSS.n578 292.5
R1968 VSS.n582 VSS.n580 292.5
R1969 VSS.n572 VSS.n571 292.5
R1970 VSS.n5721 VSS.n572 292.5
R1971 VSS.n5731 VSS.n5730 292.5
R1972 VSS.n5732 VSS.n5731 292.5
R1973 VSS.n561 VSS.n559 292.5
R1974 VSS.n563 VSS.n561 292.5
R1975 VSS.n553 VSS.n552 292.5
R1976 VSS.n5744 VSS.n553 292.5
R1977 VSS.n5754 VSS.n5753 292.5
R1978 VSS.n5755 VSS.n5754 292.5
R1979 VSS.n542 VSS.n540 292.5
R1980 VSS.n544 VSS.n542 292.5
R1981 VSS.n534 VSS.n533 292.5
R1982 VSS.n5767 VSS.n534 292.5
R1983 VSS.n5777 VSS.n5776 292.5
R1984 VSS.n5778 VSS.n5777 292.5
R1985 VSS.n523 VSS.n521 292.5
R1986 VSS.n525 VSS.n523 292.5
R1987 VSS.n5606 VSS.n5605 292.5
R1988 VSS.n5606 VSS.n5594 292.5
R1989 VSS.n1362 VSS.n1361 292.5
R1990 VSS.n5649 VSS.n1362 292.5
R1991 VSS.n5652 VSS.n5651 292.5
R1992 VSS.n5651 VSS.n5650 292.5
R1993 VSS.n5653 VSS.n1360 292.5
R1994 VSS.n1360 VSS.n1359 292.5
R1995 VSS.n5655 VSS.n5654 292.5
R1996 VSS.n5656 VSS.n5655 292.5
R1997 VSS.n1358 VSS.n1357 292.5
R1998 VSS.n5657 VSS.n1358 292.5
R1999 VSS.n5660 VSS.n5659 292.5
R2000 VSS.n5659 VSS.n5658 292.5
R2001 VSS.n5661 VSS.n1356 292.5
R2002 VSS.n1356 VSS.n1355 292.5
R2003 VSS.n5663 VSS.n5662 292.5
R2004 VSS.n5664 VSS.n5663 292.5
R2005 VSS.n1354 VSS.n1353 292.5
R2006 VSS.n5665 VSS.n1354 292.5
R2007 VSS.n5668 VSS.n5667 292.5
R2008 VSS.n5667 VSS.n5666 292.5
R2009 VSS.n5669 VSS.n1352 292.5
R2010 VSS.n1352 VSS.n1351 292.5
R2011 VSS.n5671 VSS.n5670 292.5
R2012 VSS.n5672 VSS.n5671 292.5
R2013 VSS.n1490 VSS.n1489 292.5
R2014 VSS.n1491 VSS.n1490 292.5
R2015 VSS.n1488 VSS.n1463 292.5
R2016 VSS.n1463 VSS.n1462 292.5
R2017 VSS.n1487 VSS.n1486 292.5
R2018 VSS.n1486 VSS.n1485 292.5
R2019 VSS.n1465 VSS.n1464 292.5
R2020 VSS.n1484 VSS.n1465 292.5
R2021 VSS.n1482 VSS.n1481 292.5
R2022 VSS.n1483 VSS.n1482 292.5
R2023 VSS.n1480 VSS.n1467 292.5
R2024 VSS.n1467 VSS.n1466 292.5
R2025 VSS.n1479 VSS.n1478 292.5
R2026 VSS.n1478 VSS.n1477 292.5
R2027 VSS.n1469 VSS.n1468 292.5
R2028 VSS.n1476 VSS.n1469 292.5
R2029 VSS.n1474 VSS.n1473 292.5
R2030 VSS.n1475 VSS.n1474 292.5
R2031 VSS.n1472 VSS.n1471 292.5
R2032 VSS.n1471 VSS.n1470 292.5
R2033 VSS.n1367 VSS.n1365 292.5
R2034 VSS.n1365 VSS.n1364 292.5
R2035 VSS.n5646 VSS.n5645 292.5
R2036 VSS.n5647 VSS.n5646 292.5
R2037 VSS.n1385 VSS.n1384 292.5
R2038 VSS.n5593 VSS.n1385 292.5
R2039 VSS.n1394 VSS.n1392 292.5
R2040 VSS.n5580 VSS.n1394 292.5
R2041 VSS.n5577 VSS.n5576 292.5
R2042 VSS.n5578 VSS.n5577 292.5
R2043 VSS.n1401 VSS.n1399 292.5
R2044 VSS.n5567 VSS.n1401 292.5
R2045 VSS.n5558 VSS.n5557 292.5
R2046 VSS.n5557 VSS.n5556 292.5
R2047 VSS.n1410 VSS.n1409 292.5
R2048 VSS.n1409 VSS.n1408 292.5
R2049 VSS.n5542 VSS.n5541 292.5
R2050 VSS.n5543 VSS.n5542 292.5
R2051 VSS.n1422 VSS.n1420 292.5
R2052 VSS.n5532 VSS.n1422 292.5
R2053 VSS.n5523 VSS.n5522 292.5
R2054 VSS.n5522 VSS.n5521 292.5
R2055 VSS.n1431 VSS.n1430 292.5
R2056 VSS.n1430 VSS.n1429 292.5
R2057 VSS.n5507 VSS.n5506 292.5
R2058 VSS.n5508 VSS.n5507 292.5
R2059 VSS.n1443 VSS.n1441 292.5
R2060 VSS.n5497 VSS.n1443 292.5
R2061 VSS.n5307 VSS.n5305 292.5
R2062 VSS.n5308 VSS.n5307 292.5
R2063 VSS.n5298 VSS.n5297 292.5
R2064 VSS.n5319 VSS.n5298 292.5
R2065 VSS.n5329 VSS.n5328 292.5
R2066 VSS.n5330 VSS.n5329 292.5
R2067 VSS.n5287 VSS.n5285 292.5
R2068 VSS.n5289 VSS.n5287 292.5
R2069 VSS.n5279 VSS.n5278 292.5
R2070 VSS.n5342 VSS.n5279 292.5
R2071 VSS.n5352 VSS.n5351 292.5
R2072 VSS.n5353 VSS.n5352 292.5
R2073 VSS.n5268 VSS.n5266 292.5
R2074 VSS.n5270 VSS.n5268 292.5
R2075 VSS.n5260 VSS.n5259 292.5
R2076 VSS.n5365 VSS.n5260 292.5
R2077 VSS.n5375 VSS.n5374 292.5
R2078 VSS.n5376 VSS.n5375 292.5
R2079 VSS.n5249 VSS.n5247 292.5
R2080 VSS.n5251 VSS.n5249 292.5
R2081 VSS.n5240 VSS.n5239 292.5
R2082 VSS.n5388 VSS.n5240 292.5
R2083 VSS.n5398 VSS.n5397 292.5
R2084 VSS.n5398 VSS.n5235 292.5
R2085 VSS.n1503 VSS.n1502 292.5
R2086 VSS.n5441 VSS.n1503 292.5
R2087 VSS.n5444 VSS.n5443 292.5
R2088 VSS.n5443 VSS.n5442 292.5
R2089 VSS.n5445 VSS.n1501 292.5
R2090 VSS.n1501 VSS.n1500 292.5
R2091 VSS.n5447 VSS.n5446 292.5
R2092 VSS.n5448 VSS.n5447 292.5
R2093 VSS.n1499 VSS.n1498 292.5
R2094 VSS.n5449 VSS.n1499 292.5
R2095 VSS.n5452 VSS.n5451 292.5
R2096 VSS.n5451 VSS.n5450 292.5
R2097 VSS.n5453 VSS.n1497 292.5
R2098 VSS.n1497 VSS.n1496 292.5
R2099 VSS.n5455 VSS.n5454 292.5
R2100 VSS.n5456 VSS.n5455 292.5
R2101 VSS.n1495 VSS.n1494 292.5
R2102 VSS.n5457 VSS.n1495 292.5
R2103 VSS.n5460 VSS.n5459 292.5
R2104 VSS.n5459 VSS.n5458 292.5
R2105 VSS.n5461 VSS.n1493 292.5
R2106 VSS.n1493 VSS.n1492 292.5
R2107 VSS.n5463 VSS.n5462 292.5
R2108 VSS.n5464 VSS.n5463 292.5
R2109 VSS.n1627 VSS.n1626 292.5
R2110 VSS.n1626 VSS.n1625 292.5
R2111 VSS.n1602 VSS.n1601 292.5
R2112 VSS.n1624 VSS.n1602 292.5
R2113 VSS.n1622 VSS.n1621 292.5
R2114 VSS.n1623 VSS.n1622 292.5
R2115 VSS.n1620 VSS.n1604 292.5
R2116 VSS.n1604 VSS.n1603 292.5
R2117 VSS.n1619 VSS.n1618 292.5
R2118 VSS.n1618 VSS.n1617 292.5
R2119 VSS.n1606 VSS.n1605 292.5
R2120 VSS.n1616 VSS.n1606 292.5
R2121 VSS.n1614 VSS.n1613 292.5
R2122 VSS.n1615 VSS.n1614 292.5
R2123 VSS.n1612 VSS.n1608 292.5
R2124 VSS.n1608 VSS.n1607 292.5
R2125 VSS.n1611 VSS.n1610 292.5
R2126 VSS.n1610 VSS.n1609 292.5
R2127 VSS.n1508 VSS.n1506 292.5
R2128 VSS.n1506 VSS.n1505 292.5
R2129 VSS.n5438 VSS.n5437 292.5
R2130 VSS.n5439 VSS.n5438 292.5
R2131 VSS.n1628 VSS.n1600 292.5
R2132 VSS.n1600 VSS.n1599 292.5
R2133 VSS.n1526 VSS.n1525 292.5
R2134 VSS.n5234 VSS.n1526 292.5
R2135 VSS.n1535 VSS.n1533 292.5
R2136 VSS.n5221 VSS.n1535 292.5
R2137 VSS.n5218 VSS.n5217 292.5
R2138 VSS.n5219 VSS.n5218 292.5
R2139 VSS.n1542 VSS.n1540 292.5
R2140 VSS.n5208 VSS.n1542 292.5
R2141 VSS.n5199 VSS.n5198 292.5
R2142 VSS.n5198 VSS.n5197 292.5
R2143 VSS.n1551 VSS.n1550 292.5
R2144 VSS.n1550 VSS.n1549 292.5
R2145 VSS.n5183 VSS.n5182 292.5
R2146 VSS.n5184 VSS.n5183 292.5
R2147 VSS.n1563 VSS.n1561 292.5
R2148 VSS.n5173 VSS.n1563 292.5
R2149 VSS.n5164 VSS.n5163 292.5
R2150 VSS.n5163 VSS.n5162 292.5
R2151 VSS.n1572 VSS.n1571 292.5
R2152 VSS.n1571 VSS.n1570 292.5
R2153 VSS.n5148 VSS.n5147 292.5
R2154 VSS.n5149 VSS.n5148 292.5
R2155 VSS.n1584 VSS.n1582 292.5
R2156 VSS.n5138 VSS.n1584 292.5
R2157 VSS.n1654 VSS.n1653 292.5
R2158 VSS.n3814 VSS.n3813 292.5
R2159 VSS.n3813 VSS.n3812 292.5
R2160 VSS.n3435 VSS.n3434 292.5
R2161 VSS.n3835 VSS.n3435 292.5
R2162 VSS.n3833 VSS.n3832 292.5
R2163 VSS.n3834 VSS.n3833 292.5
R2164 VSS.n3831 VSS.n3437 292.5
R2165 VSS.n3437 VSS.n3436 292.5
R2166 VSS.n3830 VSS.n3829 292.5
R2167 VSS.n3829 VSS.n3828 292.5
R2168 VSS.n3439 VSS.n3438 292.5
R2169 VSS.n3827 VSS.n3439 292.5
R2170 VSS.n3825 VSS.n3824 292.5
R2171 VSS.n3826 VSS.n3825 292.5
R2172 VSS.n3823 VSS.n3441 292.5
R2173 VSS.n3441 VSS.n3440 292.5
R2174 VSS.n3822 VSS.n3821 292.5
R2175 VSS.n3821 VSS.n3820 292.5
R2176 VSS.n3443 VSS.n3442 292.5
R2177 VSS.n3819 VSS.n3443 292.5
R2178 VSS.n3817 VSS.n3816 292.5
R2179 VSS.n3818 VSS.n3817 292.5
R2180 VSS.n3815 VSS.n3445 292.5
R2181 VSS.n3445 VSS.n3444 292.5
R2182 VSS.n4835 VSS.n4834 292.5
R2183 VSS.n4842 VSS.n4835 292.5
R2184 VSS.n3098 VSS.n3096 292.5
R2185 VSS.n3100 VSS.n3098 292.5
R2186 VSS.n4764 VSS.n4762 292.5
R2187 VSS.n4769 VSS.n4764 292.5
R2188 VSS.n4921 VSS.n4920 292.5
R2189 VSS.n4922 VSS.n4921 292.5
R2190 VSS.n4778 VSS.n4777 292.5
R2191 VSS.n4911 VSS.n4778 292.5
R2192 VSS.n4786 VSS.n4784 292.5
R2193 VSS.n4788 VSS.n4786 292.5
R2194 VSS.n4898 VSS.n4897 292.5
R2195 VSS.n4899 VSS.n4898 292.5
R2196 VSS.n4797 VSS.n4796 292.5
R2197 VSS.n4888 VSS.n4797 292.5
R2198 VSS.n4805 VSS.n4803 292.5
R2199 VSS.n4807 VSS.n4805 292.5
R2200 VSS.n4875 VSS.n4874 292.5
R2201 VSS.n4876 VSS.n4875 292.5
R2202 VSS.n4816 VSS.n4815 292.5
R2203 VSS.n4865 VSS.n4816 292.5
R2204 VSS.n4824 VSS.n4822 292.5
R2205 VSS.n4826 VSS.n4824 292.5
R2206 VSS.n4852 VSS.n4851 292.5
R2207 VSS.n4853 VSS.n4852 292.5
R2208 VSS.n3099 VSS.n3097 292.5
R2209 VSS.n5125 VSS.n3099 292.5
R2210 VSS.n5123 VSS.n5122 292.5
R2211 VSS.n5124 VSS.n5123 292.5
R2212 VSS.n5121 VSS.n3102 292.5
R2213 VSS.n3102 VSS.n3101 292.5
R2214 VSS.n5120 VSS.n5119 292.5
R2215 VSS.n5119 VSS.n5118 292.5
R2216 VSS.n3104 VSS.n3103 292.5
R2217 VSS.n5117 VSS.n3104 292.5
R2218 VSS.n5115 VSS.n5114 292.5
R2219 VSS.n5116 VSS.n5115 292.5
R2220 VSS.n5113 VSS.n3106 292.5
R2221 VSS.n3106 VSS.n3105 292.5
R2222 VSS.n5112 VSS.n5111 292.5
R2223 VSS.n5111 VSS.n5110 292.5
R2224 VSS.n3108 VSS.n3107 292.5
R2225 VSS.n5109 VSS.n3108 292.5
R2226 VSS.n5107 VSS.n5106 292.5
R2227 VSS.n5108 VSS.n5107 292.5
R2228 VSS.n5105 VSS.n3110 292.5
R2229 VSS.n3110 VSS.n3109 292.5
R2230 VSS.n5128 VSS.n5127 292.5
R2231 VSS.n5127 VSS.n5126 292.5
R2232 VSS.n5081 VSS.n3122 292.5
R2233 VSS.n3122 VSS.n3121 292.5
R2234 VSS.n5083 VSS.n5082 292.5
R2235 VSS.n5084 VSS.n5083 292.5
R2236 VSS.n3120 VSS.n3119 292.5
R2237 VSS.n5085 VSS.n3120 292.5
R2238 VSS.n5088 VSS.n5087 292.5
R2239 VSS.n5087 VSS.n5086 292.5
R2240 VSS.n5089 VSS.n3118 292.5
R2241 VSS.n3118 VSS.n3117 292.5
R2242 VSS.n5091 VSS.n5090 292.5
R2243 VSS.n5092 VSS.n5091 292.5
R2244 VSS.n3116 VSS.n3115 292.5
R2245 VSS.n5093 VSS.n3116 292.5
R2246 VSS.n5096 VSS.n5095 292.5
R2247 VSS.n5095 VSS.n5094 292.5
R2248 VSS.n5097 VSS.n3114 292.5
R2249 VSS.n3114 VSS.n3113 292.5
R2250 VSS.n5099 VSS.n5098 292.5
R2251 VSS.n5100 VSS.n5099 292.5
R2252 VSS.n3112 VSS.n3111 292.5
R2253 VSS.n5101 VSS.n3112 292.5
R2254 VSS.n5104 VSS.n5103 292.5
R2255 VSS.n5103 VSS.n5102 292.5
R2256 VSS.n5053 VSS.n5052 292.5
R2257 VSS.n5052 VSS.n5051 292.5
R2258 VSS.n5054 VSS.n3137 292.5
R2259 VSS.n3137 VSS.n3136 292.5
R2260 VSS.n5056 VSS.n5055 292.5
R2261 VSS.n5057 VSS.n5056 292.5
R2262 VSS.n3135 VSS.n3134 292.5
R2263 VSS.n5058 VSS.n3135 292.5
R2264 VSS.n5061 VSS.n5060 292.5
R2265 VSS.n5060 VSS.n5059 292.5
R2266 VSS.n5062 VSS.n3133 292.5
R2267 VSS.n3133 VSS.n3132 292.5
R2268 VSS.n5064 VSS.n5063 292.5
R2269 VSS.n5065 VSS.n5064 292.5
R2270 VSS.n3131 VSS.n3130 292.5
R2271 VSS.n5066 VSS.n3131 292.5
R2272 VSS.n5070 VSS.n5069 292.5
R2273 VSS.n5069 VSS.n5068 292.5
R2274 VSS.n5071 VSS.n3129 292.5
R2275 VSS.n5067 VSS.n3129 292.5
R2276 VSS.n5073 VSS.n5072 292.5
R2277 VSS.n5073 VSS.n3128 292.5
R2278 VSS.n5074 VSS.n3123 292.5
R2279 VSS.n5075 VSS.n5074 292.5
R2280 VSS.n4723 VSS.n4722 292.5
R2281 VSS.n4935 VSS.n4723 292.5
R2282 VSS.n4945 VSS.n4944 292.5
R2283 VSS.n4946 VSS.n4945 292.5
R2284 VSS.n4712 VSS.n4710 292.5
R2285 VSS.n4714 VSS.n4712 292.5
R2286 VSS.n4704 VSS.n4703 292.5
R2287 VSS.n4958 VSS.n4704 292.5
R2288 VSS.n4968 VSS.n4967 292.5
R2289 VSS.n4969 VSS.n4968 292.5
R2290 VSS.n4693 VSS.n4691 292.5
R2291 VSS.n4695 VSS.n4693 292.5
R2292 VSS.n4685 VSS.n4684 292.5
R2293 VSS.n4981 VSS.n4685 292.5
R2294 VSS.n4991 VSS.n4990 292.5
R2295 VSS.n4992 VSS.n4991 292.5
R2296 VSS.n4674 VSS.n4672 292.5
R2297 VSS.n4676 VSS.n4674 292.5
R2298 VSS.n4666 VSS.n4665 292.5
R2299 VSS.n5004 VSS.n4666 292.5
R2300 VSS.n5014 VSS.n5013 292.5
R2301 VSS.n5015 VSS.n5014 292.5
R2302 VSS.n4653 VSS.n4651 292.5
R2303 VSS.n4657 VSS.n4653 292.5
R2304 VSS.n3159 VSS.n3158 292.5
R2305 VSS.n4643 VSS.n3159 292.5
R2306 VSS.n4634 VSS.n4633 292.5
R2307 VSS.n4633 VSS.n4632 292.5
R2308 VSS.n3168 VSS.n3167 292.5
R2309 VSS.n3167 VSS.n3166 292.5
R2310 VSS.n4618 VSS.n4617 292.5
R2311 VSS.n4619 VSS.n4618 292.5
R2312 VSS.n3180 VSS.n3178 292.5
R2313 VSS.n4608 VSS.n3180 292.5
R2314 VSS.n4599 VSS.n4598 292.5
R2315 VSS.n4598 VSS.n4597 292.5
R2316 VSS.n3189 VSS.n3188 292.5
R2317 VSS.n3188 VSS.n3187 292.5
R2318 VSS.n4583 VSS.n4582 292.5
R2319 VSS.n4584 VSS.n4583 292.5
R2320 VSS.n3201 VSS.n3199 292.5
R2321 VSS.n4573 VSS.n3201 292.5
R2322 VSS.n4564 VSS.n4563 292.5
R2323 VSS.n4563 VSS.n4562 292.5
R2324 VSS.n3210 VSS.n3209 292.5
R2325 VSS.n3209 VSS.n3208 292.5
R2326 VSS.n4548 VSS.n4547 292.5
R2327 VSS.n4549 VSS.n4548 292.5
R2328 VSS.n3276 VSS.n3275 292.5
R2329 VSS.n3277 VSS.n3276 292.5
R2330 VSS.n3274 VSS.n3244 292.5
R2331 VSS.n3244 VSS.n3243 292.5
R2332 VSS.n3273 VSS.n3272 292.5
R2333 VSS.n3272 VSS.n3271 292.5
R2334 VSS.n3246 VSS.n3245 292.5
R2335 VSS.n3270 VSS.n3246 292.5
R2336 VSS.n3268 VSS.n3267 292.5
R2337 VSS.n3269 VSS.n3268 292.5
R2338 VSS.n3266 VSS.n3248 292.5
R2339 VSS.n3248 VSS.n3247 292.5
R2340 VSS.n3265 VSS.n3264 292.5
R2341 VSS.n3264 VSS.n3263 292.5
R2342 VSS.n3250 VSS.n3249 292.5
R2343 VSS.n3262 VSS.n3250 292.5
R2344 VSS.n3260 VSS.n3259 292.5
R2345 VSS.n3261 VSS.n3260 292.5
R2346 VSS.n3258 VSS.n3252 292.5
R2347 VSS.n3252 VSS.n3251 292.5
R2348 VSS.n3257 VSS.n3256 292.5
R2349 VSS.n3256 VSS.n3255 292.5
R2350 VSS.n3254 VSS.n3253 292.5
R2351 VSS.n3254 VSS.n3140 292.5
R2352 VSS.n3289 VSS.n3288 292.5
R2353 VSS.n4479 VSS.n3289 292.5
R2354 VSS.n4482 VSS.n4481 292.5
R2355 VSS.n4481 VSS.n4480 292.5
R2356 VSS.n4483 VSS.n3287 292.5
R2357 VSS.n3287 VSS.n3286 292.5
R2358 VSS.n4485 VSS.n4484 292.5
R2359 VSS.n4486 VSS.n4485 292.5
R2360 VSS.n3285 VSS.n3284 292.5
R2361 VSS.n4487 VSS.n3285 292.5
R2362 VSS.n4490 VSS.n4489 292.5
R2363 VSS.n4489 VSS.n4488 292.5
R2364 VSS.n4491 VSS.n3283 292.5
R2365 VSS.n3283 VSS.n3282 292.5
R2366 VSS.n4493 VSS.n4492 292.5
R2367 VSS.n4494 VSS.n4493 292.5
R2368 VSS.n3281 VSS.n3280 292.5
R2369 VSS.n4495 VSS.n3281 292.5
R2370 VSS.n4498 VSS.n4497 292.5
R2371 VSS.n4497 VSS.n4496 292.5
R2372 VSS.n4499 VSS.n3279 292.5
R2373 VSS.n3279 VSS.n3278 292.5
R2374 VSS.n4501 VSS.n4500 292.5
R2375 VSS.n4502 VSS.n4501 292.5
R2376 VSS.n3226 VSS.n3224 292.5
R2377 VSS.n4533 VSS.n3226 292.5
R2378 VSS.n4243 VSS.n4242 292.5
R2379 VSS.n4244 VSS.n4243 292.5
R2380 VSS.n4234 VSS.n4232 292.5
R2381 VSS.n4236 VSS.n4234 292.5
R2382 VSS.n4226 VSS.n4225 292.5
R2383 VSS.n4256 VSS.n4226 292.5
R2384 VSS.n4266 VSS.n4265 292.5
R2385 VSS.n4267 VSS.n4266 292.5
R2386 VSS.n4215 VSS.n4213 292.5
R2387 VSS.n4217 VSS.n4215 292.5
R2388 VSS.n4207 VSS.n4206 292.5
R2389 VSS.n4279 VSS.n4207 292.5
R2390 VSS.n4289 VSS.n4288 292.5
R2391 VSS.n4290 VSS.n4289 292.5
R2392 VSS.n4196 VSS.n4194 292.5
R2393 VSS.n4198 VSS.n4196 292.5
R2394 VSS.n4188 VSS.n4187 292.5
R2395 VSS.n4302 VSS.n4188 292.5
R2396 VSS.n4312 VSS.n4311 292.5
R2397 VSS.n4313 VSS.n4312 292.5
R2398 VSS.n4174 VSS.n4172 292.5
R2399 VSS.n4179 VSS.n4174 292.5
R2400 VSS.n4133 VSS.n4132 292.5
R2401 VSS.n4326 VSS.n4133 292.5
R2402 VSS.n4336 VSS.n4335 292.5
R2403 VSS.n4337 VSS.n4336 292.5
R2404 VSS.n4122 VSS.n4120 292.5
R2405 VSS.n4124 VSS.n4122 292.5
R2406 VSS.n4114 VSS.n4113 292.5
R2407 VSS.n4349 VSS.n4114 292.5
R2408 VSS.n4359 VSS.n4358 292.5
R2409 VSS.n4360 VSS.n4359 292.5
R2410 VSS.n4103 VSS.n4101 292.5
R2411 VSS.n4105 VSS.n4103 292.5
R2412 VSS.n4095 VSS.n4094 292.5
R2413 VSS.n4372 VSS.n4095 292.5
R2414 VSS.n4382 VSS.n4381 292.5
R2415 VSS.n4383 VSS.n4382 292.5
R2416 VSS.n4084 VSS.n4082 292.5
R2417 VSS.n4086 VSS.n4084 292.5
R2418 VSS.n4076 VSS.n4075 292.5
R2419 VSS.n4395 VSS.n4076 292.5
R2420 VSS.n4405 VSS.n4404 292.5
R2421 VSS.n4406 VSS.n4405 292.5
R2422 VSS.n4065 VSS.n4061 292.5
R2423 VSS.n4067 VSS.n4065 292.5
R2424 VSS.n4450 VSS.n4449 292.5
R2425 VSS.n4451 VSS.n4450 292.5
R2426 VSS.n3304 VSS.n3303 292.5
R2427 VSS.n4452 VSS.n3304 292.5
R2428 VSS.n4455 VSS.n4454 292.5
R2429 VSS.n4454 VSS.n4453 292.5
R2430 VSS.n4456 VSS.n3302 292.5
R2431 VSS.n3302 VSS.n3301 292.5
R2432 VSS.n4458 VSS.n4457 292.5
R2433 VSS.n4459 VSS.n4458 292.5
R2434 VSS.n3300 VSS.n3299 292.5
R2435 VSS.n4460 VSS.n3300 292.5
R2436 VSS.n4463 VSS.n4462 292.5
R2437 VSS.n4462 VSS.n4461 292.5
R2438 VSS.n4464 VSS.n3298 292.5
R2439 VSS.n3298 VSS.n3297 292.5
R2440 VSS.n4467 VSS.n4466 292.5
R2441 VSS.n4468 VSS.n4467 292.5
R2442 VSS.n4465 VSS.n3296 292.5
R2443 VSS.n4469 VSS.n3296 292.5
R2444 VSS.n4471 VSS.n3295 292.5
R2445 VSS.n4471 VSS.n4470 292.5
R2446 VSS.n4473 VSS.n4472 292.5
R2447 VSS.n4472 VSS.n3290 292.5
R2448 VSS.n3919 VSS.n3405 292.5
R2449 VSS.n3920 VSS.n3919 292.5
R2450 VSS.n3918 VSS.n3917 292.5
R2451 VSS.n3918 VSS.n3887 292.5
R2452 VSS.n3916 VSS.n3888 292.5
R2453 VSS.n3891 VSS.n3888 292.5
R2454 VSS.n3915 VSS.n3914 292.5
R2455 VSS.n3914 VSS.n3913 292.5
R2456 VSS.n3890 VSS.n3889 292.5
R2457 VSS.n3912 VSS.n3890 292.5
R2458 VSS.n3910 VSS.n3909 292.5
R2459 VSS.n3911 VSS.n3910 292.5
R2460 VSS.n3908 VSS.n3893 292.5
R2461 VSS.n3893 VSS.n3892 292.5
R2462 VSS.n3907 VSS.n3906 292.5
R2463 VSS.n3906 VSS.n3905 292.5
R2464 VSS.n3895 VSS.n3894 292.5
R2465 VSS.n3904 VSS.n3895 292.5
R2466 VSS.n3902 VSS.n3901 292.5
R2467 VSS.n3903 VSS.n3902 292.5
R2468 VSS.n3900 VSS.n3899 292.5
R2469 VSS.n3899 VSS.n3896 292.5
R2470 VSS.n3898 VSS.n3307 292.5
R2471 VSS.n3898 VSS.n3897 292.5
R2472 VSS.n3325 VSS.n3324 292.5
R2473 VSS.n3324 VSS.n3323 292.5
R2474 VSS.n4052 VSS.n4051 292.5
R2475 VSS.n4053 VSS.n4052 292.5
R2476 VSS.n3336 VSS.n3334 292.5
R2477 VSS.n4042 VSS.n3336 292.5
R2478 VSS.n4033 VSS.n4032 292.5
R2479 VSS.n4032 VSS.n4031 292.5
R2480 VSS.n3345 VSS.n3344 292.5
R2481 VSS.n3344 VSS.n3343 292.5
R2482 VSS.n4017 VSS.n4016 292.5
R2483 VSS.n4018 VSS.n4017 292.5
R2484 VSS.n3357 VSS.n3355 292.5
R2485 VSS.n4007 VSS.n3357 292.5
R2486 VSS.n3998 VSS.n3997 292.5
R2487 VSS.n3997 VSS.n3996 292.5
R2488 VSS.n3366 VSS.n3365 292.5
R2489 VSS.n3365 VSS.n3364 292.5
R2490 VSS.n3982 VSS.n3981 292.5
R2491 VSS.n3983 VSS.n3982 292.5
R2492 VSS.n3378 VSS.n3376 292.5
R2493 VSS.n3972 VSS.n3378 292.5
R2494 VSS.n3963 VSS.n3962 292.5
R2495 VSS.n3962 VSS.n3961 292.5
R2496 VSS.n3389 VSS.n3387 292.5
R2497 VSS.n3387 VSS.n3386 292.5
R2498 VSS.n3639 VSS.n3638 292.5
R2499 VSS.n3640 VSS.n3639 292.5
R2500 VSS.n3622 VSS.n3620 292.5
R2501 VSS.n3624 VSS.n3622 292.5
R2502 VSS.n3614 VSS.n3613 292.5
R2503 VSS.n3652 VSS.n3614 292.5
R2504 VSS.n3662 VSS.n3661 292.5
R2505 VSS.n3663 VSS.n3662 292.5
R2506 VSS.n3603 VSS.n3601 292.5
R2507 VSS.n3605 VSS.n3603 292.5
R2508 VSS.n3595 VSS.n3594 292.5
R2509 VSS.n3675 VSS.n3595 292.5
R2510 VSS.n3685 VSS.n3684 292.5
R2511 VSS.n3686 VSS.n3685 292.5
R2512 VSS.n3584 VSS.n3582 292.5
R2513 VSS.n3586 VSS.n3584 292.5
R2514 VSS.n3576 VSS.n3575 292.5
R2515 VSS.n3698 VSS.n3576 292.5
R2516 VSS.n3708 VSS.n3707 292.5
R2517 VSS.n3709 VSS.n3708 292.5
R2518 VSS.n3562 VSS.n3560 292.5
R2519 VSS.n3567 VSS.n3562 292.5
R2520 VSS.n3866 VSS.n3418 292.5
R2521 VSS.n3418 VSS.n3417 292.5
R2522 VSS.n3868 VSS.n3867 292.5
R2523 VSS.n3869 VSS.n3868 292.5
R2524 VSS.n3416 VSS.n3415 292.5
R2525 VSS.n3870 VSS.n3416 292.5
R2526 VSS.n3873 VSS.n3872 292.5
R2527 VSS.n3872 VSS.n3871 292.5
R2528 VSS.n3874 VSS.n3414 292.5
R2529 VSS.n3414 VSS.n3413 292.5
R2530 VSS.n3876 VSS.n3875 292.5
R2531 VSS.n3877 VSS.n3876 292.5
R2532 VSS.n3412 VSS.n3411 292.5
R2533 VSS.n3878 VSS.n3412 292.5
R2534 VSS.n3881 VSS.n3880 292.5
R2535 VSS.n3880 VSS.n3879 292.5
R2536 VSS.n3882 VSS.n3410 292.5
R2537 VSS.n3410 VSS.n3409 292.5
R2538 VSS.n3884 VSS.n3883 292.5
R2539 VSS.n3885 VSS.n3884 292.5
R2540 VSS.n3407 VSS.n3406 292.5
R2541 VSS.n3886 VSS.n3407 292.5
R2542 VSS.n3924 VSS.n3923 292.5
R2543 VSS.n3923 VSS.n3922 292.5
R2544 VSS.n3839 VSS.n3433 292.5
R2545 VSS.n3433 VSS.n3432 292.5
R2546 VSS.n3841 VSS.n3840 292.5
R2547 VSS.n3842 VSS.n3841 292.5
R2548 VSS.n3431 VSS.n3430 292.5
R2549 VSS.n3843 VSS.n3431 292.5
R2550 VSS.n3846 VSS.n3845 292.5
R2551 VSS.n3845 VSS.n3844 292.5
R2552 VSS.n3847 VSS.n3429 292.5
R2553 VSS.n3429 VSS.n3428 292.5
R2554 VSS.n3849 VSS.n3848 292.5
R2555 VSS.n3850 VSS.n3849 292.5
R2556 VSS.n3427 VSS.n3426 292.5
R2557 VSS.n3851 VSS.n3427 292.5
R2558 VSS.n3855 VSS.n3854 292.5
R2559 VSS.n3854 VSS.n3853 292.5
R2560 VSS.n3856 VSS.n3425 292.5
R2561 VSS.n3852 VSS.n3425 292.5
R2562 VSS.n3858 VSS.n3857 292.5
R2563 VSS.n3858 VSS.n3424 292.5
R2564 VSS.n3859 VSS.n3419 292.5
R2565 VSS.n3860 VSS.n3859 292.5
R2566 VSS.n3838 VSS.n3837 292.5
R2567 VSS.n3837 VSS.n3836 292.5
R2568 VSS.n3521 VSS.n3520 292.5
R2569 VSS.n3722 VSS.n3521 292.5
R2570 VSS.n3732 VSS.n3731 292.5
R2571 VSS.n3733 VSS.n3732 292.5
R2572 VSS.n3510 VSS.n3508 292.5
R2573 VSS.n3512 VSS.n3510 292.5
R2574 VSS.n3502 VSS.n3501 292.5
R2575 VSS.n3745 VSS.n3502 292.5
R2576 VSS.n3755 VSS.n3754 292.5
R2577 VSS.n3756 VSS.n3755 292.5
R2578 VSS.n3491 VSS.n3489 292.5
R2579 VSS.n3493 VSS.n3491 292.5
R2580 VSS.n3483 VSS.n3482 292.5
R2581 VSS.n3768 VSS.n3483 292.5
R2582 VSS.n3778 VSS.n3777 292.5
R2583 VSS.n3779 VSS.n3778 292.5
R2584 VSS.n3472 VSS.n3470 292.5
R2585 VSS.n3474 VSS.n3472 292.5
R2586 VSS.n3464 VSS.n3463 292.5
R2587 VSS.n3791 VSS.n3464 292.5
R2588 VSS.n3801 VSS.n3800 292.5
R2589 VSS.n3802 VSS.n3801 292.5
R2590 VSS.n3807 VSS.n3450 292.5
R2591 VSS.n3450 VSS.n3449 292.5
R2592 VSS.n3448 VSS.n3446 292.5
R2593 VSS.n17851 VSS.n17809 292.5
R2594 VSS.n17852 VSS.n17851 292.5
R2595 VSS.n17831 VSS.n17830 292.5
R2596 VSS.n17830 VSS.n17829 292.5
R2597 VSS.n17832 VSS.n17819 292.5
R2598 VSS.n17819 VSS.n17818 292.5
R2599 VSS.n17834 VSS.n17833 292.5
R2600 VSS.n17835 VSS.n17834 292.5
R2601 VSS.n17817 VSS.n17816 292.5
R2602 VSS.n17836 VSS.n17817 292.5
R2603 VSS.n17839 VSS.n17838 292.5
R2604 VSS.n17838 VSS.n17837 292.5
R2605 VSS.n17840 VSS.n17815 292.5
R2606 VSS.n17815 VSS.n17814 292.5
R2607 VSS.n17842 VSS.n17841 292.5
R2608 VSS.n17843 VSS.n17842 292.5
R2609 VSS.n17812 VSS.n17811 292.5
R2610 VSS.n17844 VSS.n17812 292.5
R2611 VSS.n17847 VSS.n17846 292.5
R2612 VSS.n17846 VSS.n17845 292.5
R2613 VSS.n17848 VSS.n17810 292.5
R2614 VSS.n17813 VSS.n17810 292.5
R2615 VSS.n17850 VSS.n17849 292.5
R2616 VSS.n17850 VSS.n17808 292.5
R2617 VSS.n17856 VSS.n17855 292.5
R2618 VSS.n17855 VSS.n17854 292.5
R2619 VSS.n17794 VSS.n17793 292.5
R2620 VSS.n17877 VSS.n17794 292.5
R2621 VSS.n17875 VSS.n17874 292.5
R2622 VSS.n17876 VSS.n17875 292.5
R2623 VSS.n17873 VSS.n17796 292.5
R2624 VSS.n17796 VSS.n17795 292.5
R2625 VSS.n17872 VSS.n17871 292.5
R2626 VSS.n17871 VSS.n17870 292.5
R2627 VSS.n17798 VSS.n17797 292.5
R2628 VSS.n17869 VSS.n17798 292.5
R2629 VSS.n17867 VSS.n17866 292.5
R2630 VSS.n17868 VSS.n17867 292.5
R2631 VSS.n17865 VSS.n17800 292.5
R2632 VSS.n17800 VSS.n17799 292.5
R2633 VSS.n17864 VSS.n17863 292.5
R2634 VSS.n17863 VSS.n17862 292.5
R2635 VSS.n17802 VSS.n17801 292.5
R2636 VSS.n17861 VSS.n17802 292.5
R2637 VSS.n17859 VSS.n17858 292.5
R2638 VSS.n17860 VSS.n17859 292.5
R2639 VSS.n17857 VSS.n17804 292.5
R2640 VSS.n17804 VSS.n17803 292.5
R2641 VSS.n17807 VSS.n17805 292.5
R2642 VSS.n17880 VSS.n17879 292.5
R2643 VSS.n17879 VSS.n17878 292.5
R2644 VSS.n17883 VSS.n17882 292.5
R2645 VSS.n17884 VSS.n17883 292.5
R2646 VSS.n17790 VSS.n17789 292.5
R2647 VSS.n17885 VSS.n17790 292.5
R2648 VSS.n17888 VSS.n17887 292.5
R2649 VSS.n17887 VSS.n17886 292.5
R2650 VSS.n17889 VSS.n17788 292.5
R2651 VSS.n17788 VSS.n17787 292.5
R2652 VSS.n17891 VSS.n17890 292.5
R2653 VSS.n17892 VSS.n17891 292.5
R2654 VSS.n17786 VSS.n17785 292.5
R2655 VSS.n17893 VSS.n17786 292.5
R2656 VSS.n17896 VSS.n17895 292.5
R2657 VSS.n17895 VSS.n17894 292.5
R2658 VSS.n17897 VSS.n17784 292.5
R2659 VSS.n17784 VSS.n17783 292.5
R2660 VSS.n17899 VSS.n17898 292.5
R2661 VSS.n17900 VSS.n17899 292.5
R2662 VSS.n17782 VSS.n17781 292.5
R2663 VSS.n17901 VSS.n17782 292.5
R2664 VSS.n17904 VSS.n17903 292.5
R2665 VSS.n17903 VSS.n17902 292.5
R2666 VSS.n17881 VSS.n17792 292.5
R2667 VSS.n17792 VSS.n17791 292.5
R2668 VSS.n17826 VSS.n17825 292.5
R2669 VSS.n17827 VSS.n17826 292.5
R2670 VSS.n17824 VSS.n17823 292.5
R2671 VSS.n17823 VSS.n17822 292.5
R2672 VSS.n17772 VSS.n17770 292.5
R2673 VSS.n17774 VSS.n17772 292.5
R2674 VSS.n17920 VSS.n17919 292.5
R2675 VSS.n17919 VSS.n17918 292.5
R2676 VSS.n17773 VSS.n17771 292.5
R2677 VSS.n17917 VSS.n17773 292.5
R2678 VSS.n17915 VSS.n17914 292.5
R2679 VSS.n17916 VSS.n17915 292.5
R2680 VSS.n17913 VSS.n17776 292.5
R2681 VSS.n17776 VSS.n17775 292.5
R2682 VSS.n17912 VSS.n17911 292.5
R2683 VSS.n17911 VSS.n17910 292.5
R2684 VSS.n17778 VSS.n17777 292.5
R2685 VSS.n17909 VSS.n17778 292.5
R2686 VSS.n17907 VSS.n17906 292.5
R2687 VSS.n17908 VSS.n17907 292.5
R2688 VSS.n17905 VSS.n17780 292.5
R2689 VSS.n17780 VSS.n17779 292.5
R2690 VSS.n17821 VSS.n17820 292.5
R2691 VSS.n17828 VSS.n17821 292.5
R2692 VSS.n16386 VSS.n16385 287.581
R2693 VSS.n16400 VSS.n16399 287.581
R2694 VSS.n16414 VSS.n16413 287.581
R2695 VSS.n16428 VSS.n16427 287.581
R2696 VSS.n16442 VSS.n16441 287.581
R2697 VSS.n16460 VSS.n16459 287.581
R2698 VSS.n16478 VSS.n16477 287.581
R2699 VSS.n16492 VSS.n16491 287.581
R2700 VSS.n16506 VSS.n16505 287.581
R2701 VSS.n16520 VSS.n16519 287.581
R2702 VSS.n16581 VSS.n16580 287.581
R2703 VSS.n16130 VSS.n16129 287.581
R2704 VSS.n16144 VSS.n16143 287.581
R2705 VSS.n16158 VSS.n16157 287.581
R2706 VSS.n16172 VSS.n16171 287.581
R2707 VSS.n16186 VSS.n16185 287.581
R2708 VSS.n16204 VSS.n16203 287.581
R2709 VSS.n16222 VSS.n16221 287.581
R2710 VSS.n16236 VSS.n16235 287.581
R2711 VSS.n16250 VSS.n16249 287.581
R2712 VSS.n16264 VSS.n16263 287.581
R2713 VSS.n16282 VSS.n16280 287.581
R2714 VSS.n16282 VSS.n16281 287.581
R2715 VSS.n15886 VSS.n15885 287.581
R2716 VSS.n15900 VSS.n15899 287.581
R2717 VSS.n15914 VSS.n15913 287.581
R2718 VSS.n15928 VSS.n15927 287.581
R2719 VSS.n15942 VSS.n15941 287.581
R2720 VSS.n15960 VSS.n15959 287.581
R2721 VSS.n15978 VSS.n15977 287.581
R2722 VSS.n15992 VSS.n15991 287.581
R2723 VSS.n16006 VSS.n16005 287.581
R2724 VSS.n16020 VSS.n16019 287.581
R2725 VSS.n16038 VSS.n16036 287.581
R2726 VSS.n16038 VSS.n16037 287.581
R2727 VSS.n15642 VSS.n15641 287.581
R2728 VSS.n15656 VSS.n15655 287.581
R2729 VSS.n15670 VSS.n15669 287.581
R2730 VSS.n15684 VSS.n15683 287.581
R2731 VSS.n15698 VSS.n15697 287.581
R2732 VSS.n15716 VSS.n15715 287.581
R2733 VSS.n15734 VSS.n15733 287.581
R2734 VSS.n15748 VSS.n15747 287.581
R2735 VSS.n15762 VSS.n15761 287.581
R2736 VSS.n15776 VSS.n15775 287.581
R2737 VSS.n15794 VSS.n15792 287.581
R2738 VSS.n15794 VSS.n15793 287.581
R2739 VSS.n15398 VSS.n15397 287.581
R2740 VSS.n15412 VSS.n15411 287.581
R2741 VSS.n15426 VSS.n15425 287.581
R2742 VSS.n15440 VSS.n15439 287.581
R2743 VSS.n15454 VSS.n15453 287.581
R2744 VSS.n15472 VSS.n15471 287.581
R2745 VSS.n15490 VSS.n15489 287.581
R2746 VSS.n15504 VSS.n15503 287.581
R2747 VSS.n15518 VSS.n15517 287.581
R2748 VSS.n15532 VSS.n15531 287.581
R2749 VSS.n15550 VSS.n15548 287.581
R2750 VSS.n15550 VSS.n15549 287.581
R2751 VSS.n15154 VSS.n15153 287.581
R2752 VSS.n15168 VSS.n15167 287.581
R2753 VSS.n15182 VSS.n15181 287.581
R2754 VSS.n15196 VSS.n15195 287.581
R2755 VSS.n15210 VSS.n15209 287.581
R2756 VSS.n15228 VSS.n15227 287.581
R2757 VSS.n15246 VSS.n15245 287.581
R2758 VSS.n15260 VSS.n15259 287.581
R2759 VSS.n15274 VSS.n15273 287.581
R2760 VSS.n15288 VSS.n15287 287.581
R2761 VSS.n15306 VSS.n15304 287.581
R2762 VSS.n15306 VSS.n15305 287.581
R2763 VSS.n14910 VSS.n14909 287.581
R2764 VSS.n14924 VSS.n14923 287.581
R2765 VSS.n14938 VSS.n14937 287.581
R2766 VSS.n14952 VSS.n14951 287.581
R2767 VSS.n14966 VSS.n14965 287.581
R2768 VSS.n14984 VSS.n14983 287.581
R2769 VSS.n15002 VSS.n15001 287.581
R2770 VSS.n15016 VSS.n15015 287.581
R2771 VSS.n15030 VSS.n15029 287.581
R2772 VSS.n15044 VSS.n15043 287.581
R2773 VSS.n15062 VSS.n15060 287.581
R2774 VSS.n15062 VSS.n15061 287.581
R2775 VSS.n14654 VSS.n14653 287.581
R2776 VSS.n14668 VSS.n14667 287.581
R2777 VSS.n14682 VSS.n14681 287.581
R2778 VSS.n14696 VSS.n14695 287.581
R2779 VSS.n14710 VSS.n14709 287.581
R2780 VSS.n14728 VSS.n14727 287.581
R2781 VSS.n14746 VSS.n14745 287.581
R2782 VSS.n14760 VSS.n14759 287.581
R2783 VSS.n14774 VSS.n14773 287.581
R2784 VSS.n14788 VSS.n14787 287.581
R2785 VSS.n14806 VSS.n14804 287.581
R2786 VSS.n14806 VSS.n14805 287.581
R2787 VSS.n12435 VSS.n12434 287.581
R2788 VSS.n12449 VSS.n12448 287.581
R2789 VSS.n12463 VSS.n12462 287.581
R2790 VSS.n12477 VSS.n12476 287.581
R2791 VSS.n12491 VSS.n12490 287.581
R2792 VSS.n12509 VSS.n12508 287.581
R2793 VSS.n12527 VSS.n12526 287.581
R2794 VSS.n12541 VSS.n12540 287.581
R2795 VSS.n12555 VSS.n12554 287.581
R2796 VSS.n12569 VSS.n12568 287.581
R2797 VSS.n12630 VSS.n12629 287.581
R2798 VSS.n12179 VSS.n12178 287.581
R2799 VSS.n12193 VSS.n12192 287.581
R2800 VSS.n12207 VSS.n12206 287.581
R2801 VSS.n12221 VSS.n12220 287.581
R2802 VSS.n12235 VSS.n12234 287.581
R2803 VSS.n12253 VSS.n12252 287.581
R2804 VSS.n12271 VSS.n12270 287.581
R2805 VSS.n12285 VSS.n12284 287.581
R2806 VSS.n12299 VSS.n12298 287.581
R2807 VSS.n12313 VSS.n12312 287.581
R2808 VSS.n12331 VSS.n12329 287.581
R2809 VSS.n12331 VSS.n12330 287.581
R2810 VSS.n11935 VSS.n11934 287.581
R2811 VSS.n11949 VSS.n11948 287.581
R2812 VSS.n11963 VSS.n11962 287.581
R2813 VSS.n11977 VSS.n11976 287.581
R2814 VSS.n11991 VSS.n11990 287.581
R2815 VSS.n12009 VSS.n12008 287.581
R2816 VSS.n12027 VSS.n12026 287.581
R2817 VSS.n12041 VSS.n12040 287.581
R2818 VSS.n12055 VSS.n12054 287.581
R2819 VSS.n12069 VSS.n12068 287.581
R2820 VSS.n12087 VSS.n12085 287.581
R2821 VSS.n12087 VSS.n12086 287.581
R2822 VSS.n11691 VSS.n11690 287.581
R2823 VSS.n11705 VSS.n11704 287.581
R2824 VSS.n11719 VSS.n11718 287.581
R2825 VSS.n11733 VSS.n11732 287.581
R2826 VSS.n11747 VSS.n11746 287.581
R2827 VSS.n11765 VSS.n11764 287.581
R2828 VSS.n11783 VSS.n11782 287.581
R2829 VSS.n11797 VSS.n11796 287.581
R2830 VSS.n11811 VSS.n11810 287.581
R2831 VSS.n11825 VSS.n11824 287.581
R2832 VSS.n11843 VSS.n11841 287.581
R2833 VSS.n11843 VSS.n11842 287.581
R2834 VSS.n11447 VSS.n11446 287.581
R2835 VSS.n11461 VSS.n11460 287.581
R2836 VSS.n11475 VSS.n11474 287.581
R2837 VSS.n11489 VSS.n11488 287.581
R2838 VSS.n11503 VSS.n11502 287.581
R2839 VSS.n11521 VSS.n11520 287.581
R2840 VSS.n11539 VSS.n11538 287.581
R2841 VSS.n11553 VSS.n11552 287.581
R2842 VSS.n11567 VSS.n11566 287.581
R2843 VSS.n11581 VSS.n11580 287.581
R2844 VSS.n11599 VSS.n11597 287.581
R2845 VSS.n11599 VSS.n11598 287.581
R2846 VSS.n11203 VSS.n11202 287.581
R2847 VSS.n11217 VSS.n11216 287.581
R2848 VSS.n11231 VSS.n11230 287.581
R2849 VSS.n11245 VSS.n11244 287.581
R2850 VSS.n11259 VSS.n11258 287.581
R2851 VSS.n11277 VSS.n11276 287.581
R2852 VSS.n11295 VSS.n11294 287.581
R2853 VSS.n11309 VSS.n11308 287.581
R2854 VSS.n11323 VSS.n11322 287.581
R2855 VSS.n11337 VSS.n11336 287.581
R2856 VSS.n11355 VSS.n11353 287.581
R2857 VSS.n11355 VSS.n11354 287.581
R2858 VSS.n10959 VSS.n10958 287.581
R2859 VSS.n10973 VSS.n10972 287.581
R2860 VSS.n10987 VSS.n10986 287.581
R2861 VSS.n11001 VSS.n11000 287.581
R2862 VSS.n11015 VSS.n11014 287.581
R2863 VSS.n11033 VSS.n11032 287.581
R2864 VSS.n11051 VSS.n11050 287.581
R2865 VSS.n11065 VSS.n11064 287.581
R2866 VSS.n11079 VSS.n11078 287.581
R2867 VSS.n11093 VSS.n11092 287.581
R2868 VSS.n11111 VSS.n11109 287.581
R2869 VSS.n11111 VSS.n11110 287.581
R2870 VSS.n10703 VSS.n10702 287.581
R2871 VSS.n10717 VSS.n10716 287.581
R2872 VSS.n10731 VSS.n10730 287.581
R2873 VSS.n10745 VSS.n10744 287.581
R2874 VSS.n10759 VSS.n10758 287.581
R2875 VSS.n10777 VSS.n10776 287.581
R2876 VSS.n10795 VSS.n10794 287.581
R2877 VSS.n10809 VSS.n10808 287.581
R2878 VSS.n10823 VSS.n10822 287.581
R2879 VSS.n10837 VSS.n10836 287.581
R2880 VSS.n10855 VSS.n10853 287.581
R2881 VSS.n10855 VSS.n10854 287.581
R2882 VSS.n9003 VSS.n9002 287.581
R2883 VSS.n9017 VSS.n9016 287.581
R2884 VSS.n9031 VSS.n9030 287.581
R2885 VSS.n9045 VSS.n9044 287.581
R2886 VSS.n9059 VSS.n9058 287.581
R2887 VSS.n9077 VSS.n9076 287.581
R2888 VSS.n9095 VSS.n9094 287.581
R2889 VSS.n9109 VSS.n9108 287.581
R2890 VSS.n9123 VSS.n9122 287.581
R2891 VSS.n9137 VSS.n9136 287.581
R2892 VSS.n9198 VSS.n9197 287.581
R2893 VSS.n8747 VSS.n8746 287.581
R2894 VSS.n8761 VSS.n8760 287.581
R2895 VSS.n8775 VSS.n8774 287.581
R2896 VSS.n8789 VSS.n8788 287.581
R2897 VSS.n8803 VSS.n8802 287.581
R2898 VSS.n8821 VSS.n8820 287.581
R2899 VSS.n8839 VSS.n8838 287.581
R2900 VSS.n8853 VSS.n8852 287.581
R2901 VSS.n8867 VSS.n8866 287.581
R2902 VSS.n8881 VSS.n8880 287.581
R2903 VSS.n8899 VSS.n8897 287.581
R2904 VSS.n8899 VSS.n8898 287.581
R2905 VSS.n8503 VSS.n8502 287.581
R2906 VSS.n8517 VSS.n8516 287.581
R2907 VSS.n8531 VSS.n8530 287.581
R2908 VSS.n8545 VSS.n8544 287.581
R2909 VSS.n8559 VSS.n8558 287.581
R2910 VSS.n8577 VSS.n8576 287.581
R2911 VSS.n8595 VSS.n8594 287.581
R2912 VSS.n8609 VSS.n8608 287.581
R2913 VSS.n8623 VSS.n8622 287.581
R2914 VSS.n8637 VSS.n8636 287.581
R2915 VSS.n8655 VSS.n8653 287.581
R2916 VSS.n8655 VSS.n8654 287.581
R2917 VSS.n8259 VSS.n8258 287.581
R2918 VSS.n8273 VSS.n8272 287.581
R2919 VSS.n8287 VSS.n8286 287.581
R2920 VSS.n8301 VSS.n8300 287.581
R2921 VSS.n8315 VSS.n8314 287.581
R2922 VSS.n8333 VSS.n8332 287.581
R2923 VSS.n8351 VSS.n8350 287.581
R2924 VSS.n8365 VSS.n8364 287.581
R2925 VSS.n8379 VSS.n8378 287.581
R2926 VSS.n8393 VSS.n8392 287.581
R2927 VSS.n8411 VSS.n8409 287.581
R2928 VSS.n8411 VSS.n8410 287.581
R2929 VSS.n8015 VSS.n8014 287.581
R2930 VSS.n8029 VSS.n8028 287.581
R2931 VSS.n8043 VSS.n8042 287.581
R2932 VSS.n8057 VSS.n8056 287.581
R2933 VSS.n8071 VSS.n8070 287.581
R2934 VSS.n8089 VSS.n8088 287.581
R2935 VSS.n8107 VSS.n8106 287.581
R2936 VSS.n8121 VSS.n8120 287.581
R2937 VSS.n8135 VSS.n8134 287.581
R2938 VSS.n8149 VSS.n8148 287.581
R2939 VSS.n8167 VSS.n8165 287.581
R2940 VSS.n8167 VSS.n8166 287.581
R2941 VSS.n7771 VSS.n7770 287.581
R2942 VSS.n7785 VSS.n7784 287.581
R2943 VSS.n7799 VSS.n7798 287.581
R2944 VSS.n7813 VSS.n7812 287.581
R2945 VSS.n7827 VSS.n7826 287.581
R2946 VSS.n7845 VSS.n7844 287.581
R2947 VSS.n7863 VSS.n7862 287.581
R2948 VSS.n7877 VSS.n7876 287.581
R2949 VSS.n7891 VSS.n7890 287.581
R2950 VSS.n7905 VSS.n7904 287.581
R2951 VSS.n7923 VSS.n7921 287.581
R2952 VSS.n7923 VSS.n7922 287.581
R2953 VSS.n7527 VSS.n7526 287.581
R2954 VSS.n7541 VSS.n7540 287.581
R2955 VSS.n7555 VSS.n7554 287.581
R2956 VSS.n7569 VSS.n7568 287.581
R2957 VSS.n7583 VSS.n7582 287.581
R2958 VSS.n7601 VSS.n7600 287.581
R2959 VSS.n7619 VSS.n7618 287.581
R2960 VSS.n7633 VSS.n7632 287.581
R2961 VSS.n7647 VSS.n7646 287.581
R2962 VSS.n7661 VSS.n7660 287.581
R2963 VSS.n7679 VSS.n7677 287.581
R2964 VSS.n7679 VSS.n7678 287.581
R2965 VSS.n7271 VSS.n7270 287.581
R2966 VSS.n7285 VSS.n7284 287.581
R2967 VSS.n7299 VSS.n7298 287.581
R2968 VSS.n7313 VSS.n7312 287.581
R2969 VSS.n7327 VSS.n7326 287.581
R2970 VSS.n7345 VSS.n7344 287.581
R2971 VSS.n7363 VSS.n7362 287.581
R2972 VSS.n7377 VSS.n7376 287.581
R2973 VSS.n7391 VSS.n7390 287.581
R2974 VSS.n7405 VSS.n7404 287.581
R2975 VSS.n7423 VSS.n7421 287.581
R2976 VSS.n7423 VSS.n7422 287.581
R2977 VSS.n1257 VSS.n1025 287.581
R2978 VSS.n1255 VSS.n1026 287.581
R2979 VSS.n1244 VSS.n1243 287.581
R2980 VSS.n1234 VSS.n1044 287.581
R2981 VSS.n1232 VSS.n1045 287.581
R2982 VSS.n1221 VSS.n1220 287.581
R2983 VSS.n1211 VSS.n1063 287.581
R2984 VSS.n1209 VSS.n1064 287.581
R2985 VSS.n1198 VSS.n1197 287.581
R2986 VSS.n1188 VSS.n1082 287.581
R2987 VSS.n1186 VSS.n1083 287.581
R2988 VSS.n1175 VSS.n1174 287.581
R2989 VSS.n919 VSS.n709 287.581
R2990 VSS.n931 VSS.n930 287.581
R2991 VSS.n942 VSS.n941 287.581
R2992 VSS.n952 VSS.n694 287.581
R2993 VSS.n954 VSS.n688 287.581
R2994 VSS.n966 VSS.n965 287.581
R2995 VSS.n977 VSS.n976 287.581
R2996 VSS.n987 VSS.n673 287.581
R2997 VSS.n989 VSS.n667 287.581
R2998 VSS.n1001 VSS.n1000 287.581
R2999 VSS.n1012 VSS.n1011 287.581
R3000 VSS.n1268 VSS.n653 287.581
R3001 VSS.n1269 VSS.n1268 287.581
R3002 VSS.n784 VSS.n783 287.581
R3003 VSS.n795 VSS.n794 287.581
R3004 VSS.n805 VSS.n766 287.581
R3005 VSS.n807 VSS.n760 287.581
R3006 VSS.n819 VSS.n818 287.581
R3007 VSS.n830 VSS.n829 287.581
R3008 VSS.n840 VSS.n745 287.581
R3009 VSS.n842 VSS.n739 287.581
R3010 VSS.n854 VSS.n853 287.581
R3011 VSS.n865 VSS.n864 287.581
R3012 VSS.n875 VSS.n723 287.581
R3013 VSS.n877 VSS.n715 287.581
R3014 VSS.n917 VSS.n715 287.581
R3015 VSS.n5596 VSS.n5594 287.581
R3016 VSS.n5780 VSS.n525 287.581
R3017 VSS.n5778 VSS.n526 287.581
R3018 VSS.n5767 VSS.n5766 287.581
R3019 VSS.n5757 VSS.n544 287.581
R3020 VSS.n5755 VSS.n545 287.581
R3021 VSS.n5744 VSS.n5743 287.581
R3022 VSS.n5734 VSS.n563 287.581
R3023 VSS.n5732 VSS.n564 287.581
R3024 VSS.n5721 VSS.n5720 287.581
R3025 VSS.n5711 VSS.n582 287.581
R3026 VSS.n5709 VSS.n583 287.581
R3027 VSS.n594 VSS.n583 287.581
R3028 VSS.n5498 VSS.n5497 287.581
R3029 VSS.n5509 VSS.n5508 287.581
R3030 VSS.n5519 VSS.n1429 287.581
R3031 VSS.n5521 VSS.n1423 287.581
R3032 VSS.n5533 VSS.n5532 287.581
R3033 VSS.n5544 VSS.n5543 287.581
R3034 VSS.n5554 VSS.n1408 287.581
R3035 VSS.n5556 VSS.n1402 287.581
R3036 VSS.n5568 VSS.n5567 287.581
R3037 VSS.n5579 VSS.n5578 287.581
R3038 VSS.n5580 VSS.n1387 287.581
R3039 VSS.n5610 VSS.n5593 287.581
R3040 VSS.n5610 VSS.n5609 287.581
R3041 VSS.n5241 VSS.n5235 287.581
R3042 VSS.n5388 VSS.n5387 287.581
R3043 VSS.n5378 VSS.n5251 287.581
R3044 VSS.n5376 VSS.n5252 287.581
R3045 VSS.n5365 VSS.n5364 287.581
R3046 VSS.n5355 VSS.n5270 287.581
R3047 VSS.n5353 VSS.n5271 287.581
R3048 VSS.n5342 VSS.n5341 287.581
R3049 VSS.n5332 VSS.n5289 287.581
R3050 VSS.n5330 VSS.n5290 287.581
R3051 VSS.n5319 VSS.n5318 287.581
R3052 VSS.n5309 VSS.n5308 287.581
R3053 VSS.n5309 VSS.n1444 287.581
R3054 VSS.n5139 VSS.n5138 287.581
R3055 VSS.n5150 VSS.n5149 287.581
R3056 VSS.n5160 VSS.n1570 287.581
R3057 VSS.n5162 VSS.n1564 287.581
R3058 VSS.n5174 VSS.n5173 287.581
R3059 VSS.n5185 VSS.n5184 287.581
R3060 VSS.n5195 VSS.n1549 287.581
R3061 VSS.n5197 VSS.n1543 287.581
R3062 VSS.n5209 VSS.n5208 287.581
R3063 VSS.n5220 VSS.n5219 287.581
R3064 VSS.n5221 VSS.n1528 287.581
R3065 VSS.n5402 VSS.n5234 287.581
R3066 VSS.n5402 VSS.n5401 287.581
R3067 VSS.n4924 VSS.n4769 287.581
R3068 VSS.n4922 VSS.n4770 287.581
R3069 VSS.n4911 VSS.n4910 287.581
R3070 VSS.n4901 VSS.n4788 287.581
R3071 VSS.n4899 VSS.n4789 287.581
R3072 VSS.n4888 VSS.n4887 287.581
R3073 VSS.n4878 VSS.n4807 287.581
R3074 VSS.n4876 VSS.n4808 287.581
R3075 VSS.n4865 VSS.n4864 287.581
R3076 VSS.n4855 VSS.n4826 287.581
R3077 VSS.n4853 VSS.n4827 287.581
R3078 VSS.n4842 VSS.n4841 287.581
R3079 VSS.n5017 VSS.n4657 287.581
R3080 VSS.n5015 VSS.n4658 287.581
R3081 VSS.n5004 VSS.n5003 287.581
R3082 VSS.n4994 VSS.n4676 287.581
R3083 VSS.n4992 VSS.n4677 287.581
R3084 VSS.n4981 VSS.n4980 287.581
R3085 VSS.n4971 VSS.n4695 287.581
R3086 VSS.n4969 VSS.n4696 287.581
R3087 VSS.n4958 VSS.n4957 287.581
R3088 VSS.n4948 VSS.n4714 287.581
R3089 VSS.n4946 VSS.n4715 287.581
R3090 VSS.n4935 VSS.n4934 287.581
R3091 VSS.n4934 VSS.n4724 287.581
R3092 VSS.n4550 VSS.n4549 287.581
R3093 VSS.n4560 VSS.n3208 287.581
R3094 VSS.n4562 VSS.n3202 287.581
R3095 VSS.n4574 VSS.n4573 287.581
R3096 VSS.n4585 VSS.n4584 287.581
R3097 VSS.n4595 VSS.n3187 287.581
R3098 VSS.n4597 VSS.n3181 287.581
R3099 VSS.n4609 VSS.n4608 287.581
R3100 VSS.n4620 VSS.n4619 287.581
R3101 VSS.n4630 VSS.n3166 287.581
R3102 VSS.n4632 VSS.n3160 287.581
R3103 VSS.n4644 VSS.n4643 287.581
R3104 VSS.n4644 VSS.n3153 287.581
R3105 VSS.n4315 VSS.n4179 287.581
R3106 VSS.n4313 VSS.n4180 287.581
R3107 VSS.n4302 VSS.n4301 287.581
R3108 VSS.n4292 VSS.n4198 287.581
R3109 VSS.n4290 VSS.n4199 287.581
R3110 VSS.n4279 VSS.n4278 287.581
R3111 VSS.n4269 VSS.n4217 287.581
R3112 VSS.n4267 VSS.n4218 287.581
R3113 VSS.n4256 VSS.n4255 287.581
R3114 VSS.n4246 VSS.n4236 287.581
R3115 VSS.n4244 VSS.n3227 287.581
R3116 VSS.n4533 VSS.n4532 287.581
R3117 VSS.n4532 VSS.n3228 287.581
R3118 VSS.n4408 VSS.n4067 287.581
R3119 VSS.n4406 VSS.n4068 287.581
R3120 VSS.n4395 VSS.n4394 287.581
R3121 VSS.n4385 VSS.n4086 287.581
R3122 VSS.n4383 VSS.n4087 287.581
R3123 VSS.n4372 VSS.n4371 287.581
R3124 VSS.n4362 VSS.n4105 287.581
R3125 VSS.n4360 VSS.n4106 287.581
R3126 VSS.n4349 VSS.n4348 287.581
R3127 VSS.n4339 VSS.n4124 287.581
R3128 VSS.n4337 VSS.n4125 287.581
R3129 VSS.n4326 VSS.n4325 287.581
R3130 VSS.n4325 VSS.n4134 287.581
R3131 VSS.n3961 VSS.n3379 287.581
R3132 VSS.n3973 VSS.n3972 287.581
R3133 VSS.n3984 VSS.n3983 287.581
R3134 VSS.n3994 VSS.n3364 287.581
R3135 VSS.n3996 VSS.n3358 287.581
R3136 VSS.n4008 VSS.n4007 287.581
R3137 VSS.n4019 VSS.n4018 287.581
R3138 VSS.n4029 VSS.n3343 287.581
R3139 VSS.n4031 VSS.n3337 287.581
R3140 VSS.n4043 VSS.n4042 287.581
R3141 VSS.n4054 VSS.n4053 287.581
R3142 VSS.n4419 VSS.n3323 287.581
R3143 VSS.n4420 VSS.n4419 287.581
R3144 VSS.n3711 VSS.n3567 287.581
R3145 VSS.n3709 VSS.n3568 287.581
R3146 VSS.n3698 VSS.n3697 287.581
R3147 VSS.n3688 VSS.n3586 287.581
R3148 VSS.n3686 VSS.n3587 287.581
R3149 VSS.n3675 VSS.n3674 287.581
R3150 VSS.n3665 VSS.n3605 287.581
R3151 VSS.n3663 VSS.n3606 287.581
R3152 VSS.n3652 VSS.n3651 287.581
R3153 VSS.n3642 VSS.n3624 287.581
R3154 VSS.n3640 VSS.n3625 287.581
R3155 VSS.n3958 VSS.n3386 287.581
R3156 VSS.n3959 VSS.n3958 287.581
R3157 VSS.n3804 VSS.n3449 287.581
R3158 VSS.n3802 VSS.n3455 287.581
R3159 VSS.n3791 VSS.n3790 287.581
R3160 VSS.n3781 VSS.n3474 287.581
R3161 VSS.n3779 VSS.n3475 287.581
R3162 VSS.n3768 VSS.n3767 287.581
R3163 VSS.n3758 VSS.n3493 287.581
R3164 VSS.n3756 VSS.n3494 287.581
R3165 VSS.n3745 VSS.n3744 287.581
R3166 VSS.n3735 VSS.n3512 287.581
R3167 VSS.n3733 VSS.n3513 287.581
R3168 VSS.n3722 VSS.n3721 287.581
R3169 VSS.n3721 VSS.n3522 287.581
R3170 VSS.n2339 VSS.n2298 258.333
R3171 VSS.n2249 VSS.n2208 258.333
R3172 VSS.n2159 VSS.n2118 258.333
R3173 VSS.n2069 VSS.n2028 258.333
R3174 VSS.n1979 VSS.n1938 258.333
R3175 VSS.n1889 VSS.n1848 258.333
R3176 VSS.n1799 VSS.n1758 258.333
R3177 VSS.n1709 VSS.n1668 258.333
R3178 VSS.n6453 VSS.n6412 258.333
R3179 VSS.n6543 VSS.n6502 258.333
R3180 VSS.n6633 VSS.n6592 258.333
R3181 VSS.n1630 VSS.n1600 257.464
R3182 VSS.n3837 VSS.n3435 257.464
R3183 VSS.n17830 VSS.n17821 257.464
R3184 VSS.n1140 VSS.n1106 251.613
R3185 VSS.n5103 VSS.n3110 251.613
R3186 VSS.n17903 VSS.n17780 251.613
R3187 VSS.n2358 VSS.n2357 249.999
R3188 VSS.n2268 VSS.n2267 249.999
R3189 VSS.n2178 VSS.n2177 249.999
R3190 VSS.n2088 VSS.n2087 249.999
R3191 VSS.n1998 VSS.n1997 249.999
R3192 VSS.n1908 VSS.n1907 249.999
R3193 VSS.n1818 VSS.n1817 249.999
R3194 VSS.n1728 VSS.n1727 249.999
R3195 VSS.n6205 VSS.n6085 249.999
R3196 VSS.n6269 VSS.n5969 249.999
R3197 VSS.n6333 VSS.n5853 249.999
R3198 VSS.n6961 VSS.n6394 249.999
R3199 VSS.n6472 VSS.n6471 249.999
R3200 VSS.n6562 VSS.n6561 249.999
R3201 VSS.n6652 VSS.n6651 249.999
R3202 VSS.n17979 VSS.n17978 221.666
R3203 VSS.n2460 VSS.n2288 205
R3204 VSS.n2550 VSS.n2198 205
R3205 VSS.n2640 VSS.n2108 205
R3206 VSS.n2730 VSS.n2018 205
R3207 VSS.n2820 VSS.n1928 205
R3208 VSS.n2910 VSS.n1838 205
R3209 VSS.n3000 VSS.n1748 205
R3210 VSS.n3090 VSS.n1658 205
R3211 VSS.n6246 VSS.n6108 205
R3212 VSS.n6310 VSS.n5992 205
R3213 VSS.n6374 VSS.n5876 205
R3214 VSS.n6994 VSS.n6993 205
R3215 VSS.n6934 VSS.n6402 205
R3216 VSS.n6844 VSS.n6492 205
R3217 VSS.n6754 VSS.n6582 205
R3218 VSS.n16385 VSS.n16384 201.307
R3219 VSS.n16399 VSS.n16398 201.307
R3220 VSS.n16413 VSS.n16412 201.307
R3221 VSS.n16427 VSS.n16426 201.307
R3222 VSS.n16441 VSS.n16440 201.307
R3223 VSS.n16459 VSS.n16458 201.307
R3224 VSS.n16455 VSS.n16454 201.307
R3225 VSS.n16477 VSS.n16476 201.307
R3226 VSS.n16491 VSS.n16490 201.307
R3227 VSS.n16505 VSS.n16504 201.307
R3228 VSS.n16519 VSS.n16518 201.307
R3229 VSS.n16580 VSS.n16579 201.307
R3230 VSS.n16129 VSS.n16128 201.307
R3231 VSS.n16143 VSS.n16142 201.307
R3232 VSS.n16157 VSS.n16156 201.307
R3233 VSS.n16171 VSS.n16170 201.307
R3234 VSS.n16185 VSS.n16184 201.307
R3235 VSS.n16203 VSS.n16202 201.307
R3236 VSS.n16199 VSS.n16198 201.307
R3237 VSS.n16221 VSS.n16220 201.307
R3238 VSS.n16235 VSS.n16234 201.307
R3239 VSS.n16249 VSS.n16248 201.307
R3240 VSS.n16263 VSS.n16262 201.307
R3241 VSS.n16280 VSS.n16279 201.307
R3242 VSS.n15885 VSS.n15884 201.307
R3243 VSS.n15899 VSS.n15898 201.307
R3244 VSS.n15913 VSS.n15912 201.307
R3245 VSS.n15927 VSS.n15926 201.307
R3246 VSS.n15941 VSS.n15940 201.307
R3247 VSS.n15959 VSS.n15958 201.307
R3248 VSS.n15955 VSS.n15954 201.307
R3249 VSS.n15977 VSS.n15976 201.307
R3250 VSS.n15991 VSS.n15990 201.307
R3251 VSS.n16005 VSS.n16004 201.307
R3252 VSS.n16019 VSS.n16018 201.307
R3253 VSS.n16036 VSS.n16035 201.307
R3254 VSS.n15641 VSS.n15640 201.307
R3255 VSS.n15655 VSS.n15654 201.307
R3256 VSS.n15669 VSS.n15668 201.307
R3257 VSS.n15683 VSS.n15682 201.307
R3258 VSS.n15697 VSS.n15696 201.307
R3259 VSS.n15715 VSS.n15714 201.307
R3260 VSS.n15711 VSS.n15710 201.307
R3261 VSS.n15733 VSS.n15732 201.307
R3262 VSS.n15747 VSS.n15746 201.307
R3263 VSS.n15761 VSS.n15760 201.307
R3264 VSS.n15775 VSS.n15774 201.307
R3265 VSS.n15792 VSS.n15791 201.307
R3266 VSS.n15397 VSS.n15396 201.307
R3267 VSS.n15411 VSS.n15410 201.307
R3268 VSS.n15425 VSS.n15424 201.307
R3269 VSS.n15439 VSS.n15438 201.307
R3270 VSS.n15453 VSS.n15452 201.307
R3271 VSS.n15471 VSS.n15470 201.307
R3272 VSS.n15467 VSS.n15466 201.307
R3273 VSS.n15489 VSS.n15488 201.307
R3274 VSS.n15503 VSS.n15502 201.307
R3275 VSS.n15517 VSS.n15516 201.307
R3276 VSS.n15531 VSS.n15530 201.307
R3277 VSS.n15548 VSS.n15547 201.307
R3278 VSS.n15153 VSS.n15152 201.307
R3279 VSS.n15167 VSS.n15166 201.307
R3280 VSS.n15181 VSS.n15180 201.307
R3281 VSS.n15195 VSS.n15194 201.307
R3282 VSS.n15209 VSS.n15208 201.307
R3283 VSS.n15227 VSS.n15226 201.307
R3284 VSS.n15223 VSS.n15222 201.307
R3285 VSS.n15245 VSS.n15244 201.307
R3286 VSS.n15259 VSS.n15258 201.307
R3287 VSS.n15273 VSS.n15272 201.307
R3288 VSS.n15287 VSS.n15286 201.307
R3289 VSS.n15304 VSS.n15303 201.307
R3290 VSS.n14909 VSS.n14908 201.307
R3291 VSS.n14923 VSS.n14922 201.307
R3292 VSS.n14937 VSS.n14936 201.307
R3293 VSS.n14951 VSS.n14950 201.307
R3294 VSS.n14965 VSS.n14964 201.307
R3295 VSS.n14983 VSS.n14982 201.307
R3296 VSS.n14979 VSS.n14978 201.307
R3297 VSS.n15001 VSS.n15000 201.307
R3298 VSS.n15015 VSS.n15014 201.307
R3299 VSS.n15029 VSS.n15028 201.307
R3300 VSS.n15043 VSS.n15042 201.307
R3301 VSS.n15060 VSS.n15059 201.307
R3302 VSS.n14653 VSS.n14652 201.307
R3303 VSS.n14667 VSS.n14666 201.307
R3304 VSS.n14681 VSS.n14680 201.307
R3305 VSS.n14695 VSS.n14694 201.307
R3306 VSS.n14709 VSS.n14708 201.307
R3307 VSS.n14727 VSS.n14726 201.307
R3308 VSS.n14723 VSS.n14722 201.307
R3309 VSS.n14745 VSS.n14744 201.307
R3310 VSS.n14759 VSS.n14758 201.307
R3311 VSS.n14773 VSS.n14772 201.307
R3312 VSS.n14787 VSS.n14786 201.307
R3313 VSS.n14804 VSS.n14803 201.307
R3314 VSS.n12434 VSS.n12433 201.307
R3315 VSS.n12448 VSS.n12447 201.307
R3316 VSS.n12462 VSS.n12461 201.307
R3317 VSS.n12476 VSS.n12475 201.307
R3318 VSS.n12490 VSS.n12489 201.307
R3319 VSS.n12508 VSS.n12507 201.307
R3320 VSS.n12504 VSS.n12503 201.307
R3321 VSS.n12526 VSS.n12525 201.307
R3322 VSS.n12540 VSS.n12539 201.307
R3323 VSS.n12554 VSS.n12553 201.307
R3324 VSS.n12568 VSS.n12567 201.307
R3325 VSS.n12629 VSS.n12628 201.307
R3326 VSS.n12178 VSS.n12177 201.307
R3327 VSS.n12192 VSS.n12191 201.307
R3328 VSS.n12206 VSS.n12205 201.307
R3329 VSS.n12220 VSS.n12219 201.307
R3330 VSS.n12234 VSS.n12233 201.307
R3331 VSS.n12252 VSS.n12251 201.307
R3332 VSS.n12248 VSS.n12247 201.307
R3333 VSS.n12270 VSS.n12269 201.307
R3334 VSS.n12284 VSS.n12283 201.307
R3335 VSS.n12298 VSS.n12297 201.307
R3336 VSS.n12312 VSS.n12311 201.307
R3337 VSS.n12329 VSS.n12328 201.307
R3338 VSS.n11934 VSS.n11933 201.307
R3339 VSS.n11948 VSS.n11947 201.307
R3340 VSS.n11962 VSS.n11961 201.307
R3341 VSS.n11976 VSS.n11975 201.307
R3342 VSS.n11990 VSS.n11989 201.307
R3343 VSS.n12008 VSS.n12007 201.307
R3344 VSS.n12004 VSS.n12003 201.307
R3345 VSS.n12026 VSS.n12025 201.307
R3346 VSS.n12040 VSS.n12039 201.307
R3347 VSS.n12054 VSS.n12053 201.307
R3348 VSS.n12068 VSS.n12067 201.307
R3349 VSS.n12085 VSS.n12084 201.307
R3350 VSS.n11690 VSS.n11689 201.307
R3351 VSS.n11704 VSS.n11703 201.307
R3352 VSS.n11718 VSS.n11717 201.307
R3353 VSS.n11732 VSS.n11731 201.307
R3354 VSS.n11746 VSS.n11745 201.307
R3355 VSS.n11764 VSS.n11763 201.307
R3356 VSS.n11760 VSS.n11759 201.307
R3357 VSS.n11782 VSS.n11781 201.307
R3358 VSS.n11796 VSS.n11795 201.307
R3359 VSS.n11810 VSS.n11809 201.307
R3360 VSS.n11824 VSS.n11823 201.307
R3361 VSS.n11841 VSS.n11840 201.307
R3362 VSS.n11446 VSS.n11445 201.307
R3363 VSS.n11460 VSS.n11459 201.307
R3364 VSS.n11474 VSS.n11473 201.307
R3365 VSS.n11488 VSS.n11487 201.307
R3366 VSS.n11502 VSS.n11501 201.307
R3367 VSS.n11520 VSS.n11519 201.307
R3368 VSS.n11516 VSS.n11515 201.307
R3369 VSS.n11538 VSS.n11537 201.307
R3370 VSS.n11552 VSS.n11551 201.307
R3371 VSS.n11566 VSS.n11565 201.307
R3372 VSS.n11580 VSS.n11579 201.307
R3373 VSS.n11597 VSS.n11596 201.307
R3374 VSS.n11202 VSS.n11201 201.307
R3375 VSS.n11216 VSS.n11215 201.307
R3376 VSS.n11230 VSS.n11229 201.307
R3377 VSS.n11244 VSS.n11243 201.307
R3378 VSS.n11258 VSS.n11257 201.307
R3379 VSS.n11276 VSS.n11275 201.307
R3380 VSS.n11272 VSS.n11271 201.307
R3381 VSS.n11294 VSS.n11293 201.307
R3382 VSS.n11308 VSS.n11307 201.307
R3383 VSS.n11322 VSS.n11321 201.307
R3384 VSS.n11336 VSS.n11335 201.307
R3385 VSS.n11353 VSS.n11352 201.307
R3386 VSS.n10958 VSS.n10957 201.307
R3387 VSS.n10972 VSS.n10971 201.307
R3388 VSS.n10986 VSS.n10985 201.307
R3389 VSS.n11000 VSS.n10999 201.307
R3390 VSS.n11014 VSS.n11013 201.307
R3391 VSS.n11032 VSS.n11031 201.307
R3392 VSS.n11028 VSS.n11027 201.307
R3393 VSS.n11050 VSS.n11049 201.307
R3394 VSS.n11064 VSS.n11063 201.307
R3395 VSS.n11078 VSS.n11077 201.307
R3396 VSS.n11092 VSS.n11091 201.307
R3397 VSS.n11109 VSS.n11108 201.307
R3398 VSS.n10702 VSS.n10701 201.307
R3399 VSS.n10716 VSS.n10715 201.307
R3400 VSS.n10730 VSS.n10729 201.307
R3401 VSS.n10744 VSS.n10743 201.307
R3402 VSS.n10758 VSS.n10757 201.307
R3403 VSS.n10776 VSS.n10775 201.307
R3404 VSS.n10772 VSS.n10771 201.307
R3405 VSS.n10794 VSS.n10793 201.307
R3406 VSS.n10808 VSS.n10807 201.307
R3407 VSS.n10822 VSS.n10821 201.307
R3408 VSS.n10836 VSS.n10835 201.307
R3409 VSS.n10853 VSS.n10852 201.307
R3410 VSS.n9002 VSS.n9001 201.307
R3411 VSS.n9016 VSS.n9015 201.307
R3412 VSS.n9030 VSS.n9029 201.307
R3413 VSS.n9044 VSS.n9043 201.307
R3414 VSS.n9058 VSS.n9057 201.307
R3415 VSS.n9076 VSS.n9075 201.307
R3416 VSS.n9072 VSS.n9071 201.307
R3417 VSS.n9094 VSS.n9093 201.307
R3418 VSS.n9108 VSS.n9107 201.307
R3419 VSS.n9122 VSS.n9121 201.307
R3420 VSS.n9136 VSS.n9135 201.307
R3421 VSS.n9197 VSS.n9196 201.307
R3422 VSS.n8746 VSS.n8745 201.307
R3423 VSS.n8760 VSS.n8759 201.307
R3424 VSS.n8774 VSS.n8773 201.307
R3425 VSS.n8788 VSS.n8787 201.307
R3426 VSS.n8802 VSS.n8801 201.307
R3427 VSS.n8820 VSS.n8819 201.307
R3428 VSS.n8816 VSS.n8815 201.307
R3429 VSS.n8838 VSS.n8837 201.307
R3430 VSS.n8852 VSS.n8851 201.307
R3431 VSS.n8866 VSS.n8865 201.307
R3432 VSS.n8880 VSS.n8879 201.307
R3433 VSS.n8897 VSS.n8896 201.307
R3434 VSS.n8502 VSS.n8501 201.307
R3435 VSS.n8516 VSS.n8515 201.307
R3436 VSS.n8530 VSS.n8529 201.307
R3437 VSS.n8544 VSS.n8543 201.307
R3438 VSS.n8558 VSS.n8557 201.307
R3439 VSS.n8576 VSS.n8575 201.307
R3440 VSS.n8572 VSS.n8571 201.307
R3441 VSS.n8594 VSS.n8593 201.307
R3442 VSS.n8608 VSS.n8607 201.307
R3443 VSS.n8622 VSS.n8621 201.307
R3444 VSS.n8636 VSS.n8635 201.307
R3445 VSS.n8653 VSS.n8652 201.307
R3446 VSS.n8258 VSS.n8257 201.307
R3447 VSS.n8272 VSS.n8271 201.307
R3448 VSS.n8286 VSS.n8285 201.307
R3449 VSS.n8300 VSS.n8299 201.307
R3450 VSS.n8314 VSS.n8313 201.307
R3451 VSS.n8332 VSS.n8331 201.307
R3452 VSS.n8328 VSS.n8327 201.307
R3453 VSS.n8350 VSS.n8349 201.307
R3454 VSS.n8364 VSS.n8363 201.307
R3455 VSS.n8378 VSS.n8377 201.307
R3456 VSS.n8392 VSS.n8391 201.307
R3457 VSS.n8409 VSS.n8408 201.307
R3458 VSS.n8014 VSS.n8013 201.307
R3459 VSS.n8028 VSS.n8027 201.307
R3460 VSS.n8042 VSS.n8041 201.307
R3461 VSS.n8056 VSS.n8055 201.307
R3462 VSS.n8070 VSS.n8069 201.307
R3463 VSS.n8088 VSS.n8087 201.307
R3464 VSS.n8084 VSS.n8083 201.307
R3465 VSS.n8106 VSS.n8105 201.307
R3466 VSS.n8120 VSS.n8119 201.307
R3467 VSS.n8134 VSS.n8133 201.307
R3468 VSS.n8148 VSS.n8147 201.307
R3469 VSS.n8165 VSS.n8164 201.307
R3470 VSS.n7770 VSS.n7769 201.307
R3471 VSS.n7784 VSS.n7783 201.307
R3472 VSS.n7798 VSS.n7797 201.307
R3473 VSS.n7812 VSS.n7811 201.307
R3474 VSS.n7826 VSS.n7825 201.307
R3475 VSS.n7844 VSS.n7843 201.307
R3476 VSS.n7840 VSS.n7839 201.307
R3477 VSS.n7862 VSS.n7861 201.307
R3478 VSS.n7876 VSS.n7875 201.307
R3479 VSS.n7890 VSS.n7889 201.307
R3480 VSS.n7904 VSS.n7903 201.307
R3481 VSS.n7921 VSS.n7920 201.307
R3482 VSS.n7526 VSS.n7525 201.307
R3483 VSS.n7540 VSS.n7539 201.307
R3484 VSS.n7554 VSS.n7553 201.307
R3485 VSS.n7568 VSS.n7567 201.307
R3486 VSS.n7582 VSS.n7581 201.307
R3487 VSS.n7600 VSS.n7599 201.307
R3488 VSS.n7596 VSS.n7595 201.307
R3489 VSS.n7618 VSS.n7617 201.307
R3490 VSS.n7632 VSS.n7631 201.307
R3491 VSS.n7646 VSS.n7645 201.307
R3492 VSS.n7660 VSS.n7659 201.307
R3493 VSS.n7677 VSS.n7676 201.307
R3494 VSS.n7270 VSS.n7269 201.307
R3495 VSS.n7284 VSS.n7283 201.307
R3496 VSS.n7298 VSS.n7297 201.307
R3497 VSS.n7312 VSS.n7311 201.307
R3498 VSS.n7326 VSS.n7325 201.307
R3499 VSS.n7344 VSS.n7343 201.307
R3500 VSS.n7340 VSS.n7339 201.307
R3501 VSS.n7362 VSS.n7361 201.307
R3502 VSS.n7376 VSS.n7375 201.307
R3503 VSS.n7390 VSS.n7389 201.307
R3504 VSS.n7404 VSS.n7403 201.307
R3505 VSS.n7421 VSS.n7420 201.307
R3506 VSS.n1025 VSS.n652 201.307
R3507 VSS.n1256 VSS.n1255 201.307
R3508 VSS.n1245 VSS.n1244 201.307
R3509 VSS.n1044 VSS.n1035 201.307
R3510 VSS.n1233 VSS.n1232 201.307
R3511 VSS.n1222 VSS.n1221 201.307
R3512 VSS.n1063 VSS.n1054 201.307
R3513 VSS.n1210 VSS.n1209 201.307
R3514 VSS.n1199 VSS.n1198 201.307
R3515 VSS.n1082 VSS.n1073 201.307
R3516 VSS.n1187 VSS.n1186 201.307
R3517 VSS.n1176 VSS.n1175 201.307
R3518 VSS.n919 VSS.n918 201.307
R3519 VSS.n930 VSS.n929 201.307
R3520 VSS.n941 VSS.n702 201.307
R3521 VSS.n943 VSS.n694 201.307
R3522 VSS.n954 VSS.n953 201.307
R3523 VSS.n965 VSS.n964 201.307
R3524 VSS.n976 VSS.n681 201.307
R3525 VSS.n978 VSS.n673 201.307
R3526 VSS.n989 VSS.n988 201.307
R3527 VSS.n1000 VSS.n999 201.307
R3528 VSS.n1011 VSS.n660 201.307
R3529 VSS.n1013 VSS.n653 201.307
R3530 VSS.n783 VSS.n782 201.307
R3531 VSS.n794 VSS.n774 201.307
R3532 VSS.n796 VSS.n766 201.307
R3533 VSS.n807 VSS.n806 201.307
R3534 VSS.n818 VSS.n817 201.307
R3535 VSS.n829 VSS.n753 201.307
R3536 VSS.n831 VSS.n745 201.307
R3537 VSS.n842 VSS.n841 201.307
R3538 VSS.n853 VSS.n852 201.307
R3539 VSS.n864 VSS.n732 201.307
R3540 VSS.n866 VSS.n723 201.307
R3541 VSS.n877 VSS.n876 201.307
R3542 VSS.n5608 VSS.n5594 201.307
R3543 VSS.n5597 VSS.n525 201.307
R3544 VSS.n5779 VSS.n5778 201.307
R3545 VSS.n5768 VSS.n5767 201.307
R3546 VSS.n544 VSS.n535 201.307
R3547 VSS.n5756 VSS.n5755 201.307
R3548 VSS.n5745 VSS.n5744 201.307
R3549 VSS.n563 VSS.n554 201.307
R3550 VSS.n5733 VSS.n5732 201.307
R3551 VSS.n5722 VSS.n5721 201.307
R3552 VSS.n582 VSS.n573 201.307
R3553 VSS.n5710 VSS.n5709 201.307
R3554 VSS.n5497 VSS.n5496 201.307
R3555 VSS.n5508 VSS.n1437 201.307
R3556 VSS.n5510 VSS.n1429 201.307
R3557 VSS.n5521 VSS.n5520 201.307
R3558 VSS.n5532 VSS.n5531 201.307
R3559 VSS.n5543 VSS.n1416 201.307
R3560 VSS.n5545 VSS.n1408 201.307
R3561 VSS.n5556 VSS.n5555 201.307
R3562 VSS.n5567 VSS.n5566 201.307
R3563 VSS.n5578 VSS.n1395 201.307
R3564 VSS.n5581 VSS.n5580 201.307
R3565 VSS.n5593 VSS.n5592 201.307
R3566 VSS.n5400 VSS.n5235 201.307
R3567 VSS.n5389 VSS.n5388 201.307
R3568 VSS.n5251 VSS.n5242 201.307
R3569 VSS.n5377 VSS.n5376 201.307
R3570 VSS.n5366 VSS.n5365 201.307
R3571 VSS.n5270 VSS.n5261 201.307
R3572 VSS.n5354 VSS.n5353 201.307
R3573 VSS.n5343 VSS.n5342 201.307
R3574 VSS.n5289 VSS.n5280 201.307
R3575 VSS.n5331 VSS.n5330 201.307
R3576 VSS.n5320 VSS.n5319 201.307
R3577 VSS.n5308 VSS.n5299 201.307
R3578 VSS.n5138 VSS.n5137 201.307
R3579 VSS.n5149 VSS.n1578 201.307
R3580 VSS.n5151 VSS.n1570 201.307
R3581 VSS.n5162 VSS.n5161 201.307
R3582 VSS.n5173 VSS.n5172 201.307
R3583 VSS.n5184 VSS.n1557 201.307
R3584 VSS.n5186 VSS.n1549 201.307
R3585 VSS.n5197 VSS.n5196 201.307
R3586 VSS.n5208 VSS.n5207 201.307
R3587 VSS.n5219 VSS.n1536 201.307
R3588 VSS.n5222 VSS.n5221 201.307
R3589 VSS.n5234 VSS.n5233 201.307
R3590 VSS.n4769 VSS.n4768 201.307
R3591 VSS.n4923 VSS.n4922 201.307
R3592 VSS.n4912 VSS.n4911 201.307
R3593 VSS.n4788 VSS.n4779 201.307
R3594 VSS.n4900 VSS.n4899 201.307
R3595 VSS.n4889 VSS.n4888 201.307
R3596 VSS.n4807 VSS.n4798 201.307
R3597 VSS.n4877 VSS.n4876 201.307
R3598 VSS.n4866 VSS.n4865 201.307
R3599 VSS.n4826 VSS.n4817 201.307
R3600 VSS.n4854 VSS.n4853 201.307
R3601 VSS.n4843 VSS.n4842 201.307
R3602 VSS.n4657 VSS.n4656 201.307
R3603 VSS.n5016 VSS.n5015 201.307
R3604 VSS.n5005 VSS.n5004 201.307
R3605 VSS.n4676 VSS.n4667 201.307
R3606 VSS.n4993 VSS.n4992 201.307
R3607 VSS.n4982 VSS.n4981 201.307
R3608 VSS.n4695 VSS.n4686 201.307
R3609 VSS.n4970 VSS.n4969 201.307
R3610 VSS.n4959 VSS.n4958 201.307
R3611 VSS.n4714 VSS.n4705 201.307
R3612 VSS.n4947 VSS.n4946 201.307
R3613 VSS.n4936 VSS.n4935 201.307
R3614 VSS.n4549 VSS.n3216 201.307
R3615 VSS.n4551 VSS.n3208 201.307
R3616 VSS.n4562 VSS.n4561 201.307
R3617 VSS.n4573 VSS.n4572 201.307
R3618 VSS.n4584 VSS.n3195 201.307
R3619 VSS.n4586 VSS.n3187 201.307
R3620 VSS.n4597 VSS.n4596 201.307
R3621 VSS.n4608 VSS.n4607 201.307
R3622 VSS.n4619 VSS.n3174 201.307
R3623 VSS.n4621 VSS.n3166 201.307
R3624 VSS.n4632 VSS.n4631 201.307
R3625 VSS.n4643 VSS.n4642 201.307
R3626 VSS.n4179 VSS.n4178 201.307
R3627 VSS.n4314 VSS.n4313 201.307
R3628 VSS.n4303 VSS.n4302 201.307
R3629 VSS.n4198 VSS.n4189 201.307
R3630 VSS.n4291 VSS.n4290 201.307
R3631 VSS.n4280 VSS.n4279 201.307
R3632 VSS.n4217 VSS.n4208 201.307
R3633 VSS.n4268 VSS.n4267 201.307
R3634 VSS.n4257 VSS.n4256 201.307
R3635 VSS.n4236 VSS.n4227 201.307
R3636 VSS.n4245 VSS.n4244 201.307
R3637 VSS.n4534 VSS.n4533 201.307
R3638 VSS.n4067 VSS.n3322 201.307
R3639 VSS.n4407 VSS.n4406 201.307
R3640 VSS.n4396 VSS.n4395 201.307
R3641 VSS.n4086 VSS.n4077 201.307
R3642 VSS.n4384 VSS.n4383 201.307
R3643 VSS.n4373 VSS.n4372 201.307
R3644 VSS.n4105 VSS.n4096 201.307
R3645 VSS.n4361 VSS.n4360 201.307
R3646 VSS.n4350 VSS.n4349 201.307
R3647 VSS.n4124 VSS.n4115 201.307
R3648 VSS.n4338 VSS.n4337 201.307
R3649 VSS.n4327 VSS.n4326 201.307
R3650 VSS.n3961 VSS.n3960 201.307
R3651 VSS.n3972 VSS.n3971 201.307
R3652 VSS.n3983 VSS.n3372 201.307
R3653 VSS.n3985 VSS.n3364 201.307
R3654 VSS.n3996 VSS.n3995 201.307
R3655 VSS.n4007 VSS.n4006 201.307
R3656 VSS.n4018 VSS.n3351 201.307
R3657 VSS.n4020 VSS.n3343 201.307
R3658 VSS.n4031 VSS.n4030 201.307
R3659 VSS.n4042 VSS.n4041 201.307
R3660 VSS.n4053 VSS.n3330 201.307
R3661 VSS.n4055 VSS.n3323 201.307
R3662 VSS.n3567 VSS.n3566 201.307
R3663 VSS.n3710 VSS.n3709 201.307
R3664 VSS.n3699 VSS.n3698 201.307
R3665 VSS.n3586 VSS.n3577 201.307
R3666 VSS.n3687 VSS.n3686 201.307
R3667 VSS.n3676 VSS.n3675 201.307
R3668 VSS.n3605 VSS.n3596 201.307
R3669 VSS.n3664 VSS.n3663 201.307
R3670 VSS.n3653 VSS.n3652 201.307
R3671 VSS.n3624 VSS.n3615 201.307
R3672 VSS.n3641 VSS.n3640 201.307
R3673 VSS.n3628 VSS.n3386 201.307
R3674 VSS.n3810 VSS.n3449 201.307
R3675 VSS.n3803 VSS.n3802 201.307
R3676 VSS.n3792 VSS.n3791 201.307
R3677 VSS.n3474 VSS.n3465 201.307
R3678 VSS.n3780 VSS.n3779 201.307
R3679 VSS.n3769 VSS.n3768 201.307
R3680 VSS.n3493 VSS.n3484 201.307
R3681 VSS.n3757 VSS.n3756 201.307
R3682 VSS.n3746 VSS.n3745 201.307
R3683 VSS.n3512 VSS.n3503 201.307
R3684 VSS.n3734 VSS.n3733 201.307
R3685 VSS.n3723 VSS.n3722 201.307
R3686 VSS.n17855 VSS.n17806 195.049
R3687 VSS.n17879 VSS.n17794 187.247
R3688 VSS.t24 VSS.n2308 185
R3689 VSS.n2400 VSS.n2399 185
R3690 VSS.n2397 VSS.n2312 185
R3691 VSS.n2405 VSS.n2403 185
R3692 VSS.n2394 VSS.n2393 185
R3693 VSS.n2390 VSS.n2389 185
R3694 VSS.n2387 VSS.n2386 185
R3695 VSS.n2447 VSS.n2446 185
R3696 VSS.n2456 VSS.n2455 185
R3697 VSS.n2377 VSS.n2376 185
R3698 VSS.t24 VSS.n2309 185
R3699 VSS.n2458 VSS.n2306 185
R3700 VSS.t24 VSS.n2306 185
R3701 VSS.t24 VSS.n2310 185
R3702 VSS.n2458 VSS.n2310 185
R3703 VSS.n2458 VSS.n2305 185
R3704 VSS.t24 VSS.n2305 185
R3705 VSS.t24 VSS.n2311 185
R3706 VSS.n2458 VSS.n2311 185
R3707 VSS.n2458 VSS.n2304 185
R3708 VSS.t24 VSS.n2304 185
R3709 VSS.t24 VSS.n2459 185
R3710 VSS.n2459 VSS.n2458 185
R3711 VSS.n2458 VSS.n2308 185
R3712 VSS.t26 VSS.n2218 185
R3713 VSS.n2490 VSS.n2489 185
R3714 VSS.n2487 VSS.n2222 185
R3715 VSS.n2495 VSS.n2493 185
R3716 VSS.n2484 VSS.n2483 185
R3717 VSS.n2480 VSS.n2479 185
R3718 VSS.n2477 VSS.n2476 185
R3719 VSS.n2537 VSS.n2536 185
R3720 VSS.n2546 VSS.n2545 185
R3721 VSS.n2467 VSS.n2466 185
R3722 VSS.t26 VSS.n2219 185
R3723 VSS.n2548 VSS.n2216 185
R3724 VSS.t26 VSS.n2216 185
R3725 VSS.t26 VSS.n2220 185
R3726 VSS.n2548 VSS.n2220 185
R3727 VSS.n2548 VSS.n2215 185
R3728 VSS.t26 VSS.n2215 185
R3729 VSS.t26 VSS.n2221 185
R3730 VSS.n2548 VSS.n2221 185
R3731 VSS.n2548 VSS.n2214 185
R3732 VSS.t26 VSS.n2214 185
R3733 VSS.t26 VSS.n2549 185
R3734 VSS.n2549 VSS.n2548 185
R3735 VSS.n2548 VSS.n2218 185
R3736 VSS.t22 VSS.n2128 185
R3737 VSS.n2580 VSS.n2579 185
R3738 VSS.n2577 VSS.n2132 185
R3739 VSS.n2585 VSS.n2583 185
R3740 VSS.n2574 VSS.n2573 185
R3741 VSS.n2570 VSS.n2569 185
R3742 VSS.n2567 VSS.n2566 185
R3743 VSS.n2627 VSS.n2626 185
R3744 VSS.n2636 VSS.n2635 185
R3745 VSS.n2557 VSS.n2556 185
R3746 VSS.t22 VSS.n2129 185
R3747 VSS.n2638 VSS.n2126 185
R3748 VSS.t22 VSS.n2126 185
R3749 VSS.t22 VSS.n2130 185
R3750 VSS.n2638 VSS.n2130 185
R3751 VSS.n2638 VSS.n2125 185
R3752 VSS.t22 VSS.n2125 185
R3753 VSS.t22 VSS.n2131 185
R3754 VSS.n2638 VSS.n2131 185
R3755 VSS.n2638 VSS.n2124 185
R3756 VSS.t22 VSS.n2124 185
R3757 VSS.t22 VSS.n2639 185
R3758 VSS.n2639 VSS.n2638 185
R3759 VSS.n2638 VSS.n2128 185
R3760 VSS.t18 VSS.n2038 185
R3761 VSS.n2670 VSS.n2669 185
R3762 VSS.n2667 VSS.n2042 185
R3763 VSS.n2675 VSS.n2673 185
R3764 VSS.n2664 VSS.n2663 185
R3765 VSS.n2660 VSS.n2659 185
R3766 VSS.n2657 VSS.n2656 185
R3767 VSS.n2717 VSS.n2716 185
R3768 VSS.n2726 VSS.n2725 185
R3769 VSS.n2647 VSS.n2646 185
R3770 VSS.t18 VSS.n2039 185
R3771 VSS.n2728 VSS.n2036 185
R3772 VSS.t18 VSS.n2036 185
R3773 VSS.t18 VSS.n2040 185
R3774 VSS.n2728 VSS.n2040 185
R3775 VSS.n2728 VSS.n2035 185
R3776 VSS.t18 VSS.n2035 185
R3777 VSS.t18 VSS.n2041 185
R3778 VSS.n2728 VSS.n2041 185
R3779 VSS.n2728 VSS.n2034 185
R3780 VSS.t18 VSS.n2034 185
R3781 VSS.t18 VSS.n2729 185
R3782 VSS.n2729 VSS.n2728 185
R3783 VSS.n2728 VSS.n2038 185
R3784 VSS.t20 VSS.n1948 185
R3785 VSS.n2760 VSS.n2759 185
R3786 VSS.n2757 VSS.n1952 185
R3787 VSS.n2765 VSS.n2763 185
R3788 VSS.n2754 VSS.n2753 185
R3789 VSS.n2750 VSS.n2749 185
R3790 VSS.n2747 VSS.n2746 185
R3791 VSS.n2807 VSS.n2806 185
R3792 VSS.n2816 VSS.n2815 185
R3793 VSS.n2737 VSS.n2736 185
R3794 VSS.t20 VSS.n1949 185
R3795 VSS.n2818 VSS.n1946 185
R3796 VSS.t20 VSS.n1946 185
R3797 VSS.t20 VSS.n1950 185
R3798 VSS.n2818 VSS.n1950 185
R3799 VSS.n2818 VSS.n1945 185
R3800 VSS.t20 VSS.n1945 185
R3801 VSS.t20 VSS.n1951 185
R3802 VSS.n2818 VSS.n1951 185
R3803 VSS.n2818 VSS.n1944 185
R3804 VSS.t20 VSS.n1944 185
R3805 VSS.t20 VSS.n2819 185
R3806 VSS.n2819 VSS.n2818 185
R3807 VSS.n2818 VSS.n1948 185
R3808 VSS.t28 VSS.n1858 185
R3809 VSS.n2850 VSS.n2849 185
R3810 VSS.n2847 VSS.n1862 185
R3811 VSS.n2855 VSS.n2853 185
R3812 VSS.n2844 VSS.n2843 185
R3813 VSS.n2840 VSS.n2839 185
R3814 VSS.n2837 VSS.n2836 185
R3815 VSS.n2897 VSS.n2896 185
R3816 VSS.n2906 VSS.n2905 185
R3817 VSS.n2827 VSS.n2826 185
R3818 VSS.t28 VSS.n1859 185
R3819 VSS.n2908 VSS.n1856 185
R3820 VSS.t28 VSS.n1856 185
R3821 VSS.t28 VSS.n1860 185
R3822 VSS.n2908 VSS.n1860 185
R3823 VSS.n2908 VSS.n1855 185
R3824 VSS.t28 VSS.n1855 185
R3825 VSS.t28 VSS.n1861 185
R3826 VSS.n2908 VSS.n1861 185
R3827 VSS.n2908 VSS.n1854 185
R3828 VSS.t28 VSS.n1854 185
R3829 VSS.t28 VSS.n2909 185
R3830 VSS.n2909 VSS.n2908 185
R3831 VSS.n2908 VSS.n1858 185
R3832 VSS.t30 VSS.n1768 185
R3833 VSS.n2940 VSS.n2939 185
R3834 VSS.n2937 VSS.n1772 185
R3835 VSS.n2945 VSS.n2943 185
R3836 VSS.n2934 VSS.n2933 185
R3837 VSS.n2930 VSS.n2929 185
R3838 VSS.n2927 VSS.n2926 185
R3839 VSS.n2987 VSS.n2986 185
R3840 VSS.n2996 VSS.n2995 185
R3841 VSS.n2917 VSS.n2916 185
R3842 VSS.t30 VSS.n1769 185
R3843 VSS.n2998 VSS.n1766 185
R3844 VSS.t30 VSS.n1766 185
R3845 VSS.t30 VSS.n1770 185
R3846 VSS.n2998 VSS.n1770 185
R3847 VSS.n2998 VSS.n1765 185
R3848 VSS.t30 VSS.n1765 185
R3849 VSS.t30 VSS.n1771 185
R3850 VSS.n2998 VSS.n1771 185
R3851 VSS.n2998 VSS.n1764 185
R3852 VSS.t30 VSS.n1764 185
R3853 VSS.t30 VSS.n2999 185
R3854 VSS.n2999 VSS.n2998 185
R3855 VSS.n2998 VSS.n1768 185
R3856 VSS.t16 VSS.n1678 185
R3857 VSS.n3030 VSS.n3029 185
R3858 VSS.n3027 VSS.n1682 185
R3859 VSS.n3035 VSS.n3033 185
R3860 VSS.n3024 VSS.n3023 185
R3861 VSS.n3020 VSS.n3019 185
R3862 VSS.n3017 VSS.n3016 185
R3863 VSS.n3077 VSS.n3076 185
R3864 VSS.n3086 VSS.n3085 185
R3865 VSS.n3007 VSS.n3006 185
R3866 VSS.t16 VSS.n1679 185
R3867 VSS.n3088 VSS.n1676 185
R3868 VSS.t16 VSS.n1676 185
R3869 VSS.t16 VSS.n1680 185
R3870 VSS.n3088 VSS.n1680 185
R3871 VSS.n3088 VSS.n1675 185
R3872 VSS.t16 VSS.n1675 185
R3873 VSS.t16 VSS.n1681 185
R3874 VSS.n3088 VSS.n1681 185
R3875 VSS.n3088 VSS.n1674 185
R3876 VSS.t16 VSS.n1674 185
R3877 VSS.t16 VSS.n3089 185
R3878 VSS.n3089 VSS.n3088 185
R3879 VSS.n3088 VSS.n1678 185
R3880 VSS.n6186 VSS.n6185 185
R3881 VSS.n6170 VSS.n6169 185
R3882 VSS.n6154 VSS.n6153 185
R3883 VSS.n6138 VSS.n6137 185
R3884 VSS.n6250 VSS.n6249 185
R3885 VSS.n6130 VSS.n6129 185
R3886 VSS.n6146 VSS.n6145 185
R3887 VSS.n6162 VSS.n6161 185
R3888 VSS.n6178 VSS.n6177 185
R3889 VSS.n6070 VSS.n6069 185
R3890 VSS.n6054 VSS.n6053 185
R3891 VSS.n6038 VSS.n6037 185
R3892 VSS.n6022 VSS.n6021 185
R3893 VSS.n6314 VSS.n6313 185
R3894 VSS.n6014 VSS.n6013 185
R3895 VSS.n6030 VSS.n6029 185
R3896 VSS.n6046 VSS.n6045 185
R3897 VSS.n6062 VSS.n6061 185
R3898 VSS.n5954 VSS.n5953 185
R3899 VSS.n5938 VSS.n5937 185
R3900 VSS.n5922 VSS.n5921 185
R3901 VSS.n5906 VSS.n5905 185
R3902 VSS.n6378 VSS.n6377 185
R3903 VSS.n5898 VSS.n5897 185
R3904 VSS.n5914 VSS.n5913 185
R3905 VSS.n5930 VSS.n5929 185
R3906 VSS.n5946 VSS.n5945 185
R3907 VSS.n6998 VSS.n6997 185
R3908 VSS.n7010 VSS.n7009 185
R3909 VSS.n7022 VSS.n7021 185
R3910 VSS.n7034 VSS.n7033 185
R3911 VSS.n6942 VSS.n6940 185
R3912 VSS.n7040 VSS.n7039 185
R3913 VSS.n7028 VSS.n7027 185
R3914 VSS.n7016 VSS.n7015 185
R3915 VSS.n7004 VSS.n7003 185
R3916 VSS.t66 VSS.n6422 185
R3917 VSS.n6878 VSS.n6877 185
R3918 VSS.n6875 VSS.n6426 185
R3919 VSS.n6872 VSS.n6871 185
R3920 VSS.n6868 VSS.n6867 185
R3921 VSS.n6864 VSS.n6863 185
R3922 VSS.n6861 VSS.n6860 185
R3923 VSS.n6920 VSS.n6919 185
R3924 VSS.n6929 VSS.n6928 185
R3925 VSS.n6850 VSS.n6429 185
R3926 VSS.n6932 VSS.n6429 185
R3927 VSS.t66 VSS.n6423 185
R3928 VSS.n6932 VSS.n6423 185
R3929 VSS.n6932 VSS.n6420 185
R3930 VSS.t66 VSS.n6420 185
R3931 VSS.t66 VSS.n6424 185
R3932 VSS.n6932 VSS.n6424 185
R3933 VSS.n6932 VSS.n6419 185
R3934 VSS.t66 VSS.n6419 185
R3935 VSS.t66 VSS.n6425 185
R3936 VSS.n6932 VSS.n6425 185
R3937 VSS.n6932 VSS.n6418 185
R3938 VSS.t66 VSS.n6418 185
R3939 VSS.t66 VSS.n6933 185
R3940 VSS.n6933 VSS.n6932 185
R3941 VSS.t70 VSS.n6512 185
R3942 VSS.n6788 VSS.n6787 185
R3943 VSS.n6785 VSS.n6516 185
R3944 VSS.n6782 VSS.n6781 185
R3945 VSS.n6778 VSS.n6777 185
R3946 VSS.n6774 VSS.n6773 185
R3947 VSS.n6771 VSS.n6770 185
R3948 VSS.n6830 VSS.n6829 185
R3949 VSS.n6839 VSS.n6838 185
R3950 VSS.n6760 VSS.n6519 185
R3951 VSS.n6842 VSS.n6519 185
R3952 VSS.t70 VSS.n6513 185
R3953 VSS.n6842 VSS.n6513 185
R3954 VSS.n6842 VSS.n6510 185
R3955 VSS.t70 VSS.n6510 185
R3956 VSS.t70 VSS.n6514 185
R3957 VSS.n6842 VSS.n6514 185
R3958 VSS.n6842 VSS.n6509 185
R3959 VSS.t70 VSS.n6509 185
R3960 VSS.t70 VSS.n6515 185
R3961 VSS.n6842 VSS.n6515 185
R3962 VSS.n6842 VSS.n6508 185
R3963 VSS.t70 VSS.n6508 185
R3964 VSS.t70 VSS.n6843 185
R3965 VSS.n6843 VSS.n6842 185
R3966 VSS.t72 VSS.n6602 185
R3967 VSS.n6698 VSS.n6697 185
R3968 VSS.n6695 VSS.n6606 185
R3969 VSS.n6692 VSS.n6691 185
R3970 VSS.n6688 VSS.n6687 185
R3971 VSS.n6684 VSS.n6683 185
R3972 VSS.n6681 VSS.n6680 185
R3973 VSS.n6740 VSS.n6739 185
R3974 VSS.n6749 VSS.n6748 185
R3975 VSS.n6670 VSS.n6609 185
R3976 VSS.n6752 VSS.n6609 185
R3977 VSS.t72 VSS.n6603 185
R3978 VSS.n6752 VSS.n6603 185
R3979 VSS.n6752 VSS.n6600 185
R3980 VSS.t72 VSS.n6600 185
R3981 VSS.t72 VSS.n6604 185
R3982 VSS.n6752 VSS.n6604 185
R3983 VSS.n6752 VSS.n6599 185
R3984 VSS.t72 VSS.n6599 185
R3985 VSS.t72 VSS.n6605 185
R3986 VSS.n6752 VSS.n6605 185
R3987 VSS.n6752 VSS.n6598 185
R3988 VSS.t72 VSS.n6598 185
R3989 VSS.t72 VSS.n6753 185
R3990 VSS.n6753 VSS.n6752 185
R3991 VSS.n427 VSS.n348 185
R3992 VSS.n350 VSS.n349 185
R3993 VSS.n354 VSS.n353 185
R3994 VSS.n358 VSS.n357 185
R3995 VSS.n404 VSS.n403 185
R3996 VSS.n395 VSS.n366 185
R3997 VSS.n368 VSS.n367 185
R3998 VSS.n372 VSS.n371 185
R3999 VSS.n385 VSS.n384 185
R4000 VSS.n392 VSS.n391 185
R4001 VSS.n394 VSS.n393 185
R4002 VSS.n405 VSS.n360 185
R4003 VSS.n406 VSS.n361 185
R4004 VSS.n414 VSS.n413 185
R4005 VSS.n421 VSS.n420 185
R4006 VSS.n429 VSS.n428 185
R4007 VSS.n17948 VSS.n17925 185
R4008 VSS.n18017 VSS.n17923 185
R4009 VSS.n18017 VSS.t78 185
R4010 VSS.n18164 VSS.n18163 185
R4011 VSS.n18160 VSS.n18159 185
R4012 VSS.n18187 VSS.n18158 185
R4013 VSS.n18196 VSS.n18195 185
R4014 VSS.n18150 VSS.n18149 185
R4015 VSS.n18144 VSS.n18143 185
R4016 VSS.n18215 VSS.n18214 185
R4017 VSS.n18223 VSS.n18137 185
R4018 VSS.n18177 VSS.n18176 185
R4019 VSS.n18184 VSS.n18183 185
R4020 VSS.n18186 VSS.n18185 185
R4021 VSS.n18197 VSS.n18152 185
R4022 VSS.n18198 VSS.n18153 185
R4023 VSS.n18206 VSS.n18205 185
R4024 VSS.n18213 VSS.n18142 185
R4025 VSS.n18222 VSS.n18221 185
R4026 VSS.n14650 VSS.n14649 181.396
R4027 VSS.n10699 VSS.n10698 181.396
R4028 VSS.n7267 VSS.n7266 181.396
R4029 VSS.n5136 VSS.n1586 181.396
R4030 VSS.n3809 VSS.n3447 181.396
R4031 VSS.n1651 VSS.n1650 175.544
R4032 VSS.n1650 VSS.n1589 175.544
R4033 VSS.n1646 VSS.n1589 175.544
R4034 VSS.n1646 VSS.n1591 175.544
R4035 VSS.n1642 VSS.n1591 175.544
R4036 VSS.n1642 VSS.n1594 175.544
R4037 VSS.n1638 VSS.n1594 175.544
R4038 VSS.n1638 VSS.n1596 175.544
R4039 VSS.n1634 VSS.n1596 175.544
R4040 VSS.n1634 VSS.n1598 175.544
R4041 VSS.n1630 VSS.n1598 175.544
R4042 VSS.n5443 VSS.n1503 175.544
R4043 VSS.n5443 VSS.n1501 175.544
R4044 VSS.n5447 VSS.n1501 175.544
R4045 VSS.n5447 VSS.n1499 175.544
R4046 VSS.n5451 VSS.n1499 175.544
R4047 VSS.n5451 VSS.n1497 175.544
R4048 VSS.n5455 VSS.n1497 175.544
R4049 VSS.n5455 VSS.n1495 175.544
R4050 VSS.n5459 VSS.n1495 175.544
R4051 VSS.n5459 VSS.n1493 175.544
R4052 VSS.n5463 VSS.n1493 175.544
R4053 VSS.n1626 VSS.n1600 175.544
R4054 VSS.n1626 VSS.n1602 175.544
R4055 VSS.n1622 VSS.n1602 175.544
R4056 VSS.n1622 VSS.n1604 175.544
R4057 VSS.n1618 VSS.n1604 175.544
R4058 VSS.n1618 VSS.n1606 175.544
R4059 VSS.n1614 VSS.n1606 175.544
R4060 VSS.n1614 VSS.n1608 175.544
R4061 VSS.n1610 VSS.n1608 175.544
R4062 VSS.n1610 VSS.n1506 175.544
R4063 VSS.n5438 VSS.n1506 175.544
R4064 VSS.n5651 VSS.n1362 175.544
R4065 VSS.n5651 VSS.n1360 175.544
R4066 VSS.n5655 VSS.n1360 175.544
R4067 VSS.n5655 VSS.n1358 175.544
R4068 VSS.n5659 VSS.n1358 175.544
R4069 VSS.n5659 VSS.n1356 175.544
R4070 VSS.n5663 VSS.n1356 175.544
R4071 VSS.n5663 VSS.n1354 175.544
R4072 VSS.n5667 VSS.n1354 175.544
R4073 VSS.n5667 VSS.n1352 175.544
R4074 VSS.n5671 VSS.n1352 175.544
R4075 VSS.n1490 VSS.n1463 175.544
R4076 VSS.n1486 VSS.n1463 175.544
R4077 VSS.n1486 VSS.n1465 175.544
R4078 VSS.n1482 VSS.n1465 175.544
R4079 VSS.n1482 VSS.n1467 175.544
R4080 VSS.n1478 VSS.n1467 175.544
R4081 VSS.n1478 VSS.n1469 175.544
R4082 VSS.n1474 VSS.n1469 175.544
R4083 VSS.n1474 VSS.n1471 175.544
R4084 VSS.n1471 VSS.n1365 175.544
R4085 VSS.n5646 VSS.n1365 175.544
R4086 VSS.n1320 VSS.n1319 175.544
R4087 VSS.n1319 VSS.n625 175.544
R4088 VSS.n1315 VSS.n625 175.544
R4089 VSS.n1315 VSS.n627 175.544
R4090 VSS.n1311 VSS.n627 175.544
R4091 VSS.n1311 VSS.n630 175.544
R4092 VSS.n1307 VSS.n630 175.544
R4093 VSS.n1307 VSS.n632 175.544
R4094 VSS.n1303 VSS.n632 175.544
R4095 VSS.n1303 VSS.n634 175.544
R4096 VSS.n1299 VSS.n634 175.544
R4097 VSS.n1349 VSS.n608 175.544
R4098 VSS.n1345 VSS.n608 175.544
R4099 VSS.n1345 VSS.n610 175.544
R4100 VSS.n1341 VSS.n610 175.544
R4101 VSS.n1341 VSS.n612 175.544
R4102 VSS.n1337 VSS.n612 175.544
R4103 VSS.n1337 VSS.n614 175.544
R4104 VSS.n1333 VSS.n614 175.544
R4105 VSS.n1333 VSS.n616 175.544
R4106 VSS.n1329 VSS.n616 175.544
R4107 VSS.n1329 VSS.n618 175.544
R4108 VSS.n1164 VSS.n1096 175.544
R4109 VSS.n1160 VSS.n1096 175.544
R4110 VSS.n1160 VSS.n1098 175.544
R4111 VSS.n1156 VSS.n1098 175.544
R4112 VSS.n1156 VSS.n1100 175.544
R4113 VSS.n1152 VSS.n1100 175.544
R4114 VSS.n1152 VSS.n1102 175.544
R4115 VSS.n1148 VSS.n1102 175.544
R4116 VSS.n1148 VSS.n1104 175.544
R4117 VSS.n1144 VSS.n1104 175.544
R4118 VSS.n1144 VSS.n1106 175.544
R4119 VSS.n1120 VSS.n1118 175.544
R4120 VSS.n1120 VSS.n1116 175.544
R4121 VSS.n1124 VSS.n1116 175.544
R4122 VSS.n1124 VSS.n1114 175.544
R4123 VSS.n1128 VSS.n1114 175.544
R4124 VSS.n1128 VSS.n1112 175.544
R4125 VSS.n1132 VSS.n1112 175.544
R4126 VSS.n1132 VSS.n1110 175.544
R4127 VSS.n1136 VSS.n1110 175.544
R4128 VSS.n1136 VSS.n1108 175.544
R4129 VSS.n1140 VSS.n1108 175.544
R4130 VSS.n3813 VSS.n3445 175.544
R4131 VSS.n3817 VSS.n3445 175.544
R4132 VSS.n3817 VSS.n3443 175.544
R4133 VSS.n3821 VSS.n3443 175.544
R4134 VSS.n3821 VSS.n3441 175.544
R4135 VSS.n3825 VSS.n3441 175.544
R4136 VSS.n3825 VSS.n3439 175.544
R4137 VSS.n3829 VSS.n3439 175.544
R4138 VSS.n3829 VSS.n3437 175.544
R4139 VSS.n3833 VSS.n3437 175.544
R4140 VSS.n3833 VSS.n3435 175.544
R4141 VSS.n3868 VSS.n3418 175.544
R4142 VSS.n3868 VSS.n3416 175.544
R4143 VSS.n3872 VSS.n3416 175.544
R4144 VSS.n3872 VSS.n3414 175.544
R4145 VSS.n3876 VSS.n3414 175.544
R4146 VSS.n3876 VSS.n3412 175.544
R4147 VSS.n3880 VSS.n3412 175.544
R4148 VSS.n3880 VSS.n3410 175.544
R4149 VSS.n3884 VSS.n3410 175.544
R4150 VSS.n3884 VSS.n3407 175.544
R4151 VSS.n3923 VSS.n3407 175.544
R4152 VSS.n3837 VSS.n3433 175.544
R4153 VSS.n3841 VSS.n3433 175.544
R4154 VSS.n3841 VSS.n3431 175.544
R4155 VSS.n3845 VSS.n3431 175.544
R4156 VSS.n3845 VSS.n3429 175.544
R4157 VSS.n3849 VSS.n3429 175.544
R4158 VSS.n3849 VSS.n3427 175.544
R4159 VSS.n3854 VSS.n3427 175.544
R4160 VSS.n3854 VSS.n3425 175.544
R4161 VSS.n3858 VSS.n3425 175.544
R4162 VSS.n3859 VSS.n3858 175.544
R4163 VSS.n4450 VSS.n3304 175.544
R4164 VSS.n4454 VSS.n3304 175.544
R4165 VSS.n4454 VSS.n3302 175.544
R4166 VSS.n4458 VSS.n3302 175.544
R4167 VSS.n4458 VSS.n3300 175.544
R4168 VSS.n4462 VSS.n3300 175.544
R4169 VSS.n4462 VSS.n3298 175.544
R4170 VSS.n4467 VSS.n3298 175.544
R4171 VSS.n4467 VSS.n3296 175.544
R4172 VSS.n4471 VSS.n3296 175.544
R4173 VSS.n4472 VSS.n4471 175.544
R4174 VSS.n3919 VSS.n3918 175.544
R4175 VSS.n3918 VSS.n3888 175.544
R4176 VSS.n3914 VSS.n3888 175.544
R4177 VSS.n3914 VSS.n3890 175.544
R4178 VSS.n3910 VSS.n3890 175.544
R4179 VSS.n3910 VSS.n3893 175.544
R4180 VSS.n3906 VSS.n3893 175.544
R4181 VSS.n3906 VSS.n3895 175.544
R4182 VSS.n3902 VSS.n3895 175.544
R4183 VSS.n3902 VSS.n3899 175.544
R4184 VSS.n3899 VSS.n3898 175.544
R4185 VSS.n3276 VSS.n3244 175.544
R4186 VSS.n3272 VSS.n3244 175.544
R4187 VSS.n3272 VSS.n3246 175.544
R4188 VSS.n3268 VSS.n3246 175.544
R4189 VSS.n3268 VSS.n3248 175.544
R4190 VSS.n3264 VSS.n3248 175.544
R4191 VSS.n3264 VSS.n3250 175.544
R4192 VSS.n3260 VSS.n3250 175.544
R4193 VSS.n3260 VSS.n3252 175.544
R4194 VSS.n3256 VSS.n3252 175.544
R4195 VSS.n3256 VSS.n3254 175.544
R4196 VSS.n4481 VSS.n3289 175.544
R4197 VSS.n4481 VSS.n3287 175.544
R4198 VSS.n4485 VSS.n3287 175.544
R4199 VSS.n4485 VSS.n3285 175.544
R4200 VSS.n4489 VSS.n3285 175.544
R4201 VSS.n4489 VSS.n3283 175.544
R4202 VSS.n4493 VSS.n3283 175.544
R4203 VSS.n4493 VSS.n3281 175.544
R4204 VSS.n4497 VSS.n3281 175.544
R4205 VSS.n4497 VSS.n3279 175.544
R4206 VSS.n4501 VSS.n3279 175.544
R4207 VSS.n5052 VSS.n3137 175.544
R4208 VSS.n5056 VSS.n3137 175.544
R4209 VSS.n5056 VSS.n3135 175.544
R4210 VSS.n5060 VSS.n3135 175.544
R4211 VSS.n5060 VSS.n3133 175.544
R4212 VSS.n5064 VSS.n3133 175.544
R4213 VSS.n5064 VSS.n3131 175.544
R4214 VSS.n5069 VSS.n3131 175.544
R4215 VSS.n5069 VSS.n3129 175.544
R4216 VSS.n5073 VSS.n3129 175.544
R4217 VSS.n5074 VSS.n5073 175.544
R4218 VSS.n5083 VSS.n3122 175.544
R4219 VSS.n5083 VSS.n3120 175.544
R4220 VSS.n5087 VSS.n3120 175.544
R4221 VSS.n5087 VSS.n3118 175.544
R4222 VSS.n5091 VSS.n3118 175.544
R4223 VSS.n5091 VSS.n3116 175.544
R4224 VSS.n5095 VSS.n3116 175.544
R4225 VSS.n5095 VSS.n3114 175.544
R4226 VSS.n5099 VSS.n3114 175.544
R4227 VSS.n5099 VSS.n3112 175.544
R4228 VSS.n5103 VSS.n3112 175.544
R4229 VSS.n5127 VSS.n3099 175.544
R4230 VSS.n5123 VSS.n3099 175.544
R4231 VSS.n5123 VSS.n3102 175.544
R4232 VSS.n5119 VSS.n3102 175.544
R4233 VSS.n5119 VSS.n3104 175.544
R4234 VSS.n5115 VSS.n3104 175.544
R4235 VSS.n5115 VSS.n3106 175.544
R4236 VSS.n5111 VSS.n3106 175.544
R4237 VSS.n5111 VSS.n3108 175.544
R4238 VSS.n5107 VSS.n3108 175.544
R4239 VSS.n5107 VSS.n3110 175.544
R4240 VSS.n17883 VSS.n17792 175.544
R4241 VSS.n17883 VSS.n17790 175.544
R4242 VSS.n17887 VSS.n17790 175.544
R4243 VSS.n17887 VSS.n17788 175.544
R4244 VSS.n17891 VSS.n17788 175.544
R4245 VSS.n17891 VSS.n17786 175.544
R4246 VSS.n17895 VSS.n17786 175.544
R4247 VSS.n17895 VSS.n17784 175.544
R4248 VSS.n17899 VSS.n17784 175.544
R4249 VSS.n17899 VSS.n17782 175.544
R4250 VSS.n17903 VSS.n17782 175.544
R4251 VSS.n17826 VSS.n17821 175.544
R4252 VSS.n17826 VSS.n17823 175.544
R4253 VSS.n17823 VSS.n17772 175.544
R4254 VSS.n17919 VSS.n17772 175.544
R4255 VSS.n17919 VSS.n17773 175.544
R4256 VSS.n17915 VSS.n17773 175.544
R4257 VSS.n17915 VSS.n17776 175.544
R4258 VSS.n17911 VSS.n17776 175.544
R4259 VSS.n17911 VSS.n17778 175.544
R4260 VSS.n17907 VSS.n17778 175.544
R4261 VSS.n17907 VSS.n17780 175.544
R4262 VSS.n17851 VSS.n17850 175.544
R4263 VSS.n17850 VSS.n17810 175.544
R4264 VSS.n17846 VSS.n17810 175.544
R4265 VSS.n17846 VSS.n17812 175.544
R4266 VSS.n17842 VSS.n17812 175.544
R4267 VSS.n17842 VSS.n17815 175.544
R4268 VSS.n17838 VSS.n17815 175.544
R4269 VSS.n17838 VSS.n17817 175.544
R4270 VSS.n17834 VSS.n17817 175.544
R4271 VSS.n17834 VSS.n17819 175.544
R4272 VSS.n17830 VSS.n17819 175.544
R4273 VSS.n17855 VSS.n17804 175.544
R4274 VSS.n17859 VSS.n17804 175.544
R4275 VSS.n17859 VSS.n17802 175.544
R4276 VSS.n17863 VSS.n17802 175.544
R4277 VSS.n17863 VSS.n17800 175.544
R4278 VSS.n17867 VSS.n17800 175.544
R4279 VSS.n17867 VSS.n17798 175.544
R4280 VSS.n17871 VSS.n17798 175.544
R4281 VSS.n17871 VSS.n17796 175.544
R4282 VSS.n17875 VSS.n17796 175.544
R4283 VSS.n17875 VSS.n17794 175.544
R4284 VSS.n16582 VSS.n16578 167.742
R4285 VSS.n12631 VSS.n12627 167.742
R4286 VSS.n9199 VSS.n9195 167.742
R4287 VSS.n1173 VSS.n1093 167.742
R4288 VSS.n4840 VSS.n3098 167.742
R4289 VSS.n2376 VSS.n2290 151.666
R4290 VSS.n2466 VSS.n2200 151.666
R4291 VSS.n2556 VSS.n2110 151.666
R4292 VSS.n2646 VSS.n2020 151.666
R4293 VSS.n2736 VSS.n1930 151.666
R4294 VSS.n2826 VSS.n1840 151.666
R4295 VSS.n2916 VSS.n1750 151.666
R4296 VSS.n3006 VSS.n1660 151.666
R4297 VSS.n6249 VSS.n6076 151.666
R4298 VSS.n6313 VSS.n5960 151.666
R4299 VSS.n6377 VSS.n5844 151.666
R4300 VSS.n6944 VSS.n6942 151.666
R4301 VSS.n6429 VSS.n6404 151.666
R4302 VSS.n6519 VSS.n6494 151.666
R4303 VSS.n6609 VSS.n6584 151.666
R4304 VSS.n2372 VSS.n2290 150
R4305 VSS.n2370 VSS.n2369 150
R4306 VSS.n2366 VSS.n2365 150
R4307 VSS.n2362 VSS.n2361 150
R4308 VSS.n2354 VSS.n2353 150
R4309 VSS.n2350 VSS.n2349 150
R4310 VSS.n2346 VSS.n2345 150
R4311 VSS.n2342 VSS.n2298 150
R4312 VSS.n2460 VSS.n2289 150
R4313 VSS.n2329 VSS.n2328 150
R4314 VSS.n2333 VSS.n2332 150
R4315 VSS.n2337 VSS.n2336 150
R4316 VSS.n2282 VSS.n2200 150
R4317 VSS.n2280 VSS.n2279 150
R4318 VSS.n2276 VSS.n2275 150
R4319 VSS.n2272 VSS.n2271 150
R4320 VSS.n2264 VSS.n2263 150
R4321 VSS.n2260 VSS.n2259 150
R4322 VSS.n2256 VSS.n2255 150
R4323 VSS.n2252 VSS.n2208 150
R4324 VSS.n2550 VSS.n2199 150
R4325 VSS.n2239 VSS.n2238 150
R4326 VSS.n2243 VSS.n2242 150
R4327 VSS.n2247 VSS.n2246 150
R4328 VSS.n2192 VSS.n2110 150
R4329 VSS.n2190 VSS.n2189 150
R4330 VSS.n2186 VSS.n2185 150
R4331 VSS.n2182 VSS.n2181 150
R4332 VSS.n2174 VSS.n2173 150
R4333 VSS.n2170 VSS.n2169 150
R4334 VSS.n2166 VSS.n2165 150
R4335 VSS.n2162 VSS.n2118 150
R4336 VSS.n2640 VSS.n2109 150
R4337 VSS.n2149 VSS.n2148 150
R4338 VSS.n2153 VSS.n2152 150
R4339 VSS.n2157 VSS.n2156 150
R4340 VSS.n2102 VSS.n2020 150
R4341 VSS.n2100 VSS.n2099 150
R4342 VSS.n2096 VSS.n2095 150
R4343 VSS.n2092 VSS.n2091 150
R4344 VSS.n2084 VSS.n2083 150
R4345 VSS.n2080 VSS.n2079 150
R4346 VSS.n2076 VSS.n2075 150
R4347 VSS.n2072 VSS.n2028 150
R4348 VSS.n2730 VSS.n2019 150
R4349 VSS.n2059 VSS.n2058 150
R4350 VSS.n2063 VSS.n2062 150
R4351 VSS.n2067 VSS.n2066 150
R4352 VSS.n2012 VSS.n1930 150
R4353 VSS.n2010 VSS.n2009 150
R4354 VSS.n2006 VSS.n2005 150
R4355 VSS.n2002 VSS.n2001 150
R4356 VSS.n1994 VSS.n1993 150
R4357 VSS.n1990 VSS.n1989 150
R4358 VSS.n1986 VSS.n1985 150
R4359 VSS.n1982 VSS.n1938 150
R4360 VSS.n2820 VSS.n1929 150
R4361 VSS.n1969 VSS.n1968 150
R4362 VSS.n1973 VSS.n1972 150
R4363 VSS.n1977 VSS.n1976 150
R4364 VSS.n1922 VSS.n1840 150
R4365 VSS.n1920 VSS.n1919 150
R4366 VSS.n1916 VSS.n1915 150
R4367 VSS.n1912 VSS.n1911 150
R4368 VSS.n1904 VSS.n1903 150
R4369 VSS.n1900 VSS.n1899 150
R4370 VSS.n1896 VSS.n1895 150
R4371 VSS.n1892 VSS.n1848 150
R4372 VSS.n2910 VSS.n1839 150
R4373 VSS.n1879 VSS.n1878 150
R4374 VSS.n1883 VSS.n1882 150
R4375 VSS.n1887 VSS.n1886 150
R4376 VSS.n1832 VSS.n1750 150
R4377 VSS.n1830 VSS.n1829 150
R4378 VSS.n1826 VSS.n1825 150
R4379 VSS.n1822 VSS.n1821 150
R4380 VSS.n1814 VSS.n1813 150
R4381 VSS.n1810 VSS.n1809 150
R4382 VSS.n1806 VSS.n1805 150
R4383 VSS.n1802 VSS.n1758 150
R4384 VSS.n3000 VSS.n1749 150
R4385 VSS.n1789 VSS.n1788 150
R4386 VSS.n1793 VSS.n1792 150
R4387 VSS.n1797 VSS.n1796 150
R4388 VSS.n1742 VSS.n1660 150
R4389 VSS.n1740 VSS.n1739 150
R4390 VSS.n1736 VSS.n1735 150
R4391 VSS.n1732 VSS.n1731 150
R4392 VSS.n1724 VSS.n1723 150
R4393 VSS.n1720 VSS.n1719 150
R4394 VSS.n1716 VSS.n1715 150
R4395 VSS.n1712 VSS.n1668 150
R4396 VSS.n3090 VSS.n1659 150
R4397 VSS.n1699 VSS.n1698 150
R4398 VSS.n1703 VSS.n1702 150
R4399 VSS.n1707 VSS.n1706 150
R4400 VSS.n6192 VSS.n6191 150
R4401 VSS.n6196 VSS.n6195 150
R4402 VSS.n6200 VSS.n6199 150
R4403 VSS.n6202 VSS.n6085 150
R4404 VSS.n6209 VSS.n6208 150
R4405 VSS.n6213 VSS.n6212 150
R4406 VSS.n6217 VSS.n6216 150
R4407 VSS.n6221 VSS.n6220 150
R4408 VSS.n6237 VSS.n6236 150
R4409 VSS.n6233 VSS.n6232 150
R4410 VSS.n6229 VSS.n6228 150
R4411 VSS.n6225 VSS.n6224 150
R4412 VSS.n6256 VSS.n6255 150
R4413 VSS.n6260 VSS.n6259 150
R4414 VSS.n6264 VSS.n6263 150
R4415 VSS.n6266 VSS.n5969 150
R4416 VSS.n6273 VSS.n6272 150
R4417 VSS.n6277 VSS.n6276 150
R4418 VSS.n6281 VSS.n6280 150
R4419 VSS.n6285 VSS.n6284 150
R4420 VSS.n6301 VSS.n6300 150
R4421 VSS.n6297 VSS.n6296 150
R4422 VSS.n6293 VSS.n6292 150
R4423 VSS.n6289 VSS.n6288 150
R4424 VSS.n6320 VSS.n6319 150
R4425 VSS.n6324 VSS.n6323 150
R4426 VSS.n6328 VSS.n6327 150
R4427 VSS.n6330 VSS.n5853 150
R4428 VSS.n6337 VSS.n6336 150
R4429 VSS.n6341 VSS.n6340 150
R4430 VSS.n6345 VSS.n6344 150
R4431 VSS.n6349 VSS.n6348 150
R4432 VSS.n6365 VSS.n6364 150
R4433 VSS.n6361 VSS.n6360 150
R4434 VSS.n6357 VSS.n6356 150
R4435 VSS.n6353 VSS.n6352 150
R4436 VSS.n6948 VSS.n6398 150
R4437 VSS.n6951 VSS.n6950 150
R4438 VSS.n6955 VSS.n6954 150
R4439 VSS.n6957 VSS.n6394 150
R4440 VSS.n6965 VSS.n6963 150
R4441 VSS.n6969 VSS.n6392 150
R4442 VSS.n6973 VSS.n6971 150
R4443 VSS.n6977 VSS.n6390 150
R4444 VSS.n6991 VSS.n6384 150
R4445 VSS.n6987 VSS.n6986 150
R4446 VSS.n6984 VSS.n6387 150
R4447 VSS.n6980 VSS.n6979 150
R4448 VSS.n6486 VSS.n6404 150
R4449 VSS.n6484 VSS.n6483 150
R4450 VSS.n6480 VSS.n6479 150
R4451 VSS.n6476 VSS.n6475 150
R4452 VSS.n6468 VSS.n6467 150
R4453 VSS.n6464 VSS.n6463 150
R4454 VSS.n6460 VSS.n6459 150
R4455 VSS.n6456 VSS.n6412 150
R4456 VSS.n6934 VSS.n6403 150
R4457 VSS.n6443 VSS.n6442 150
R4458 VSS.n6447 VSS.n6446 150
R4459 VSS.n6451 VSS.n6450 150
R4460 VSS.n6576 VSS.n6494 150
R4461 VSS.n6574 VSS.n6573 150
R4462 VSS.n6570 VSS.n6569 150
R4463 VSS.n6566 VSS.n6565 150
R4464 VSS.n6558 VSS.n6557 150
R4465 VSS.n6554 VSS.n6553 150
R4466 VSS.n6550 VSS.n6549 150
R4467 VSS.n6546 VSS.n6502 150
R4468 VSS.n6844 VSS.n6493 150
R4469 VSS.n6533 VSS.n6532 150
R4470 VSS.n6537 VSS.n6536 150
R4471 VSS.n6541 VSS.n6540 150
R4472 VSS.n6666 VSS.n6584 150
R4473 VSS.n6664 VSS.n6663 150
R4474 VSS.n6660 VSS.n6659 150
R4475 VSS.n6656 VSS.n6655 150
R4476 VSS.n6648 VSS.n6647 150
R4477 VSS.n6644 VSS.n6643 150
R4478 VSS.n6640 VSS.n6639 150
R4479 VSS.n6636 VSS.n6592 150
R4480 VSS.n6754 VSS.n6583 150
R4481 VSS.n6623 VSS.n6622 150
R4482 VSS.n6627 VSS.n6626 150
R4483 VSS.n6631 VSS.n6630 150
R4484 VSS.n17995 VSS.n17994 150
R4485 VSS.n17991 VSS.n17990 150
R4486 VSS.n17987 VSS.n17986 150
R4487 VSS.n17983 VSS.n17982 150
R4488 VSS.n17975 VSS.n17974 150
R4489 VSS.n17971 VSS.n17970 150
R4490 VSS.n17967 VSS.n17966 150
R4491 VSS.n17963 VSS.n17962 150
R4492 VSS.n18015 VSS.n17947 150
R4493 VSS.n17951 VSS.n17950 150
R4494 VSS.n17955 VSS.n17954 150
R4495 VSS.n17959 VSS.n17958 150
R4496 VSS.n18011 VSS.n17946 150
R4497 VSS.n16371 VSS.n16370 146.25
R4498 VSS.n16370 VSS.n16369 146.25
R4499 VSS.n16368 VSS.n16367 146.25
R4500 VSS.n16367 VSS.n16366 146.25
R4501 VSS.n16365 VSS.n16364 146.25
R4502 VSS.n16364 VSS.n16363 146.25
R4503 VSS.n16362 VSS.n16361 146.25
R4504 VSS.n16361 VSS.n16360 146.25
R4505 VSS.n16359 VSS.n16358 146.25
R4506 VSS.n16358 VSS.n16357 146.25
R4507 VSS.n16356 VSS.n16355 146.25
R4508 VSS.n16355 VSS.n16354 146.25
R4509 VSS.n16353 VSS.n16352 146.25
R4510 VSS.n16352 VSS.n16351 146.25
R4511 VSS.n16350 VSS.n16349 146.25
R4512 VSS.n16349 VSS.n16348 146.25
R4513 VSS.n16347 VSS.n16346 146.25
R4514 VSS.n16346 VSS.n16345 146.25
R4515 VSS.n16344 VSS.n16343 146.25
R4516 VSS.n16343 VSS.n16342 146.25
R4517 VSS.n16341 VSS.n16340 146.25
R4518 VSS.n16340 VSS.n16339 146.25
R4519 VSS.n16374 VSS.n16373 146.25
R4520 VSS.n16373 VSS.n16372 146.25
R4521 VSS.n16277 VSS.n16276 146.25
R4522 VSS.n16116 VSS.n16115 146.25
R4523 VSS.n16115 VSS.n16114 146.25
R4524 VSS.n16113 VSS.n16112 146.25
R4525 VSS.n16112 VSS.n16111 146.25
R4526 VSS.n16110 VSS.n16109 146.25
R4527 VSS.n16109 VSS.n16108 146.25
R4528 VSS.n16107 VSS.n16106 146.25
R4529 VSS.n16106 VSS.n16105 146.25
R4530 VSS.n16104 VSS.n16103 146.25
R4531 VSS.n16103 VSS.n16102 146.25
R4532 VSS.n16101 VSS.n16100 146.25
R4533 VSS.n16100 VSS.n16099 146.25
R4534 VSS.n16098 VSS.n16097 146.25
R4535 VSS.n16097 VSS.n16096 146.25
R4536 VSS.n16095 VSS.n16094 146.25
R4537 VSS.n16094 VSS.n16093 146.25
R4538 VSS.n16092 VSS.n16091 146.25
R4539 VSS.n16091 VSS.n16090 146.25
R4540 VSS.n16089 VSS.n16088 146.25
R4541 VSS.n16088 VSS.n16087 146.25
R4542 VSS.n16086 VSS.n16085 146.25
R4543 VSS.n16085 VSS.n16084 146.25
R4544 VSS.n16119 VSS.n16118 146.25
R4545 VSS.n16118 VSS.n16117 146.25
R4546 VSS.n16033 VSS.n16032 146.25
R4547 VSS.n15871 VSS.n15870 146.25
R4548 VSS.n15870 VSS.n15869 146.25
R4549 VSS.n15868 VSS.n15867 146.25
R4550 VSS.n15867 VSS.n15866 146.25
R4551 VSS.n15865 VSS.n15864 146.25
R4552 VSS.n15864 VSS.n15863 146.25
R4553 VSS.n15862 VSS.n15861 146.25
R4554 VSS.n15861 VSS.n15860 146.25
R4555 VSS.n15859 VSS.n15858 146.25
R4556 VSS.n15858 VSS.n15857 146.25
R4557 VSS.n15856 VSS.n15855 146.25
R4558 VSS.n15855 VSS.n15854 146.25
R4559 VSS.n15853 VSS.n15852 146.25
R4560 VSS.n15852 VSS.n15851 146.25
R4561 VSS.n15850 VSS.n15849 146.25
R4562 VSS.n15849 VSS.n15848 146.25
R4563 VSS.n15847 VSS.n15846 146.25
R4564 VSS.n15846 VSS.n15845 146.25
R4565 VSS.n15844 VSS.n15843 146.25
R4566 VSS.n15843 VSS.n15842 146.25
R4567 VSS.n15841 VSS.n15840 146.25
R4568 VSS.n15840 VSS.n15839 146.25
R4569 VSS.n15874 VSS.n15873 146.25
R4570 VSS.n15873 VSS.n15872 146.25
R4571 VSS.n15789 VSS.n15788 146.25
R4572 VSS.n15628 VSS.n15627 146.25
R4573 VSS.n15627 VSS.n15626 146.25
R4574 VSS.n15625 VSS.n15624 146.25
R4575 VSS.n15624 VSS.n15623 146.25
R4576 VSS.n15622 VSS.n15621 146.25
R4577 VSS.n15621 VSS.n15620 146.25
R4578 VSS.n15619 VSS.n15618 146.25
R4579 VSS.n15618 VSS.n15617 146.25
R4580 VSS.n15616 VSS.n15615 146.25
R4581 VSS.n15615 VSS.n15614 146.25
R4582 VSS.n15613 VSS.n15612 146.25
R4583 VSS.n15612 VSS.n15611 146.25
R4584 VSS.n15610 VSS.n15609 146.25
R4585 VSS.n15609 VSS.n15608 146.25
R4586 VSS.n15607 VSS.n15606 146.25
R4587 VSS.n15606 VSS.n15605 146.25
R4588 VSS.n15604 VSS.n15603 146.25
R4589 VSS.n15603 VSS.n15602 146.25
R4590 VSS.n15601 VSS.n15600 146.25
R4591 VSS.n15600 VSS.n15599 146.25
R4592 VSS.n15598 VSS.n15597 146.25
R4593 VSS.n15597 VSS.n15596 146.25
R4594 VSS.n15631 VSS.n15630 146.25
R4595 VSS.n15630 VSS.n15629 146.25
R4596 VSS.n15545 VSS.n15544 146.25
R4597 VSS.n15383 VSS.n15382 146.25
R4598 VSS.n15382 VSS.n15381 146.25
R4599 VSS.n15380 VSS.n15379 146.25
R4600 VSS.n15379 VSS.n15378 146.25
R4601 VSS.n15377 VSS.n15376 146.25
R4602 VSS.n15376 VSS.n15375 146.25
R4603 VSS.n15374 VSS.n15373 146.25
R4604 VSS.n15373 VSS.n15372 146.25
R4605 VSS.n15371 VSS.n15370 146.25
R4606 VSS.n15370 VSS.n15369 146.25
R4607 VSS.n15368 VSS.n15367 146.25
R4608 VSS.n15367 VSS.n15366 146.25
R4609 VSS.n15365 VSS.n15364 146.25
R4610 VSS.n15364 VSS.n15363 146.25
R4611 VSS.n15362 VSS.n15361 146.25
R4612 VSS.n15361 VSS.n15360 146.25
R4613 VSS.n15359 VSS.n15358 146.25
R4614 VSS.n15358 VSS.n15357 146.25
R4615 VSS.n15356 VSS.n15355 146.25
R4616 VSS.n15355 VSS.n15354 146.25
R4617 VSS.n15353 VSS.n15352 146.25
R4618 VSS.n15352 VSS.n15351 146.25
R4619 VSS.n15386 VSS.n15385 146.25
R4620 VSS.n15385 VSS.n15384 146.25
R4621 VSS.n15301 VSS.n15300 146.25
R4622 VSS.n15140 VSS.n15139 146.25
R4623 VSS.n15139 VSS.n15138 146.25
R4624 VSS.n15137 VSS.n15136 146.25
R4625 VSS.n15136 VSS.n15135 146.25
R4626 VSS.n15134 VSS.n15133 146.25
R4627 VSS.n15133 VSS.n15132 146.25
R4628 VSS.n15131 VSS.n15130 146.25
R4629 VSS.n15130 VSS.n15129 146.25
R4630 VSS.n15128 VSS.n15127 146.25
R4631 VSS.n15127 VSS.n15126 146.25
R4632 VSS.n15125 VSS.n15124 146.25
R4633 VSS.n15124 VSS.n15123 146.25
R4634 VSS.n15122 VSS.n15121 146.25
R4635 VSS.n15121 VSS.n15120 146.25
R4636 VSS.n15119 VSS.n15118 146.25
R4637 VSS.n15118 VSS.n15117 146.25
R4638 VSS.n15116 VSS.n15115 146.25
R4639 VSS.n15115 VSS.n15114 146.25
R4640 VSS.n15113 VSS.n15112 146.25
R4641 VSS.n15112 VSS.n15111 146.25
R4642 VSS.n15110 VSS.n15109 146.25
R4643 VSS.n15109 VSS.n15108 146.25
R4644 VSS.n15143 VSS.n15142 146.25
R4645 VSS.n15142 VSS.n15141 146.25
R4646 VSS.n15057 VSS.n15056 146.25
R4647 VSS.n14895 VSS.n14894 146.25
R4648 VSS.n14894 VSS.n14893 146.25
R4649 VSS.n14892 VSS.n14891 146.25
R4650 VSS.n14891 VSS.n14890 146.25
R4651 VSS.n14889 VSS.n14888 146.25
R4652 VSS.n14888 VSS.n14887 146.25
R4653 VSS.n14886 VSS.n14885 146.25
R4654 VSS.n14885 VSS.n14884 146.25
R4655 VSS.n14883 VSS.n14882 146.25
R4656 VSS.n14882 VSS.n14881 146.25
R4657 VSS.n14880 VSS.n14879 146.25
R4658 VSS.n14879 VSS.n14878 146.25
R4659 VSS.n14877 VSS.n14876 146.25
R4660 VSS.n14876 VSS.n14875 146.25
R4661 VSS.n14874 VSS.n14873 146.25
R4662 VSS.n14873 VSS.n14872 146.25
R4663 VSS.n14871 VSS.n14870 146.25
R4664 VSS.n14870 VSS.n14869 146.25
R4665 VSS.n14868 VSS.n14867 146.25
R4666 VSS.n14867 VSS.n14866 146.25
R4667 VSS.n14865 VSS.n14864 146.25
R4668 VSS.n14864 VSS.n14863 146.25
R4669 VSS.n14898 VSS.n14897 146.25
R4670 VSS.n14897 VSS.n14896 146.25
R4671 VSS.n14801 VSS.n14800 146.25
R4672 VSS.n12420 VSS.n12419 146.25
R4673 VSS.n12419 VSS.n12418 146.25
R4674 VSS.n12417 VSS.n12416 146.25
R4675 VSS.n12416 VSS.n12415 146.25
R4676 VSS.n12414 VSS.n12413 146.25
R4677 VSS.n12413 VSS.n12412 146.25
R4678 VSS.n12411 VSS.n12410 146.25
R4679 VSS.n12410 VSS.n12409 146.25
R4680 VSS.n12408 VSS.n12407 146.25
R4681 VSS.n12407 VSS.n12406 146.25
R4682 VSS.n12405 VSS.n12404 146.25
R4683 VSS.n12404 VSS.n12403 146.25
R4684 VSS.n12402 VSS.n12401 146.25
R4685 VSS.n12401 VSS.n12400 146.25
R4686 VSS.n12399 VSS.n12398 146.25
R4687 VSS.n12398 VSS.n12397 146.25
R4688 VSS.n12396 VSS.n12395 146.25
R4689 VSS.n12395 VSS.n12394 146.25
R4690 VSS.n12393 VSS.n12392 146.25
R4691 VSS.n12392 VSS.n12391 146.25
R4692 VSS.n12390 VSS.n12389 146.25
R4693 VSS.n12389 VSS.n12388 146.25
R4694 VSS.n12423 VSS.n12422 146.25
R4695 VSS.n12422 VSS.n12421 146.25
R4696 VSS.n12326 VSS.n12325 146.25
R4697 VSS.n12165 VSS.n12164 146.25
R4698 VSS.n12164 VSS.n12163 146.25
R4699 VSS.n12162 VSS.n12161 146.25
R4700 VSS.n12161 VSS.n12160 146.25
R4701 VSS.n12159 VSS.n12158 146.25
R4702 VSS.n12158 VSS.n12157 146.25
R4703 VSS.n12156 VSS.n12155 146.25
R4704 VSS.n12155 VSS.n12154 146.25
R4705 VSS.n12153 VSS.n12152 146.25
R4706 VSS.n12152 VSS.n12151 146.25
R4707 VSS.n12150 VSS.n12149 146.25
R4708 VSS.n12149 VSS.n12148 146.25
R4709 VSS.n12147 VSS.n12146 146.25
R4710 VSS.n12146 VSS.n12145 146.25
R4711 VSS.n12144 VSS.n12143 146.25
R4712 VSS.n12143 VSS.n12142 146.25
R4713 VSS.n12141 VSS.n12140 146.25
R4714 VSS.n12140 VSS.n12139 146.25
R4715 VSS.n12138 VSS.n12137 146.25
R4716 VSS.n12137 VSS.n12136 146.25
R4717 VSS.n12135 VSS.n12134 146.25
R4718 VSS.n12134 VSS.n12133 146.25
R4719 VSS.n12168 VSS.n12167 146.25
R4720 VSS.n12167 VSS.n12166 146.25
R4721 VSS.n12082 VSS.n12081 146.25
R4722 VSS.n11920 VSS.n11919 146.25
R4723 VSS.n11919 VSS.n11918 146.25
R4724 VSS.n11917 VSS.n11916 146.25
R4725 VSS.n11916 VSS.n11915 146.25
R4726 VSS.n11914 VSS.n11913 146.25
R4727 VSS.n11913 VSS.n11912 146.25
R4728 VSS.n11911 VSS.n11910 146.25
R4729 VSS.n11910 VSS.n11909 146.25
R4730 VSS.n11908 VSS.n11907 146.25
R4731 VSS.n11907 VSS.n11906 146.25
R4732 VSS.n11905 VSS.n11904 146.25
R4733 VSS.n11904 VSS.n11903 146.25
R4734 VSS.n11902 VSS.n11901 146.25
R4735 VSS.n11901 VSS.n11900 146.25
R4736 VSS.n11899 VSS.n11898 146.25
R4737 VSS.n11898 VSS.n11897 146.25
R4738 VSS.n11896 VSS.n11895 146.25
R4739 VSS.n11895 VSS.n11894 146.25
R4740 VSS.n11893 VSS.n11892 146.25
R4741 VSS.n11892 VSS.n11891 146.25
R4742 VSS.n11890 VSS.n11889 146.25
R4743 VSS.n11889 VSS.n11888 146.25
R4744 VSS.n11923 VSS.n11922 146.25
R4745 VSS.n11922 VSS.n11921 146.25
R4746 VSS.n11838 VSS.n11837 146.25
R4747 VSS.n11677 VSS.n11676 146.25
R4748 VSS.n11676 VSS.n11675 146.25
R4749 VSS.n11674 VSS.n11673 146.25
R4750 VSS.n11673 VSS.n11672 146.25
R4751 VSS.n11671 VSS.n11670 146.25
R4752 VSS.n11670 VSS.n11669 146.25
R4753 VSS.n11668 VSS.n11667 146.25
R4754 VSS.n11667 VSS.n11666 146.25
R4755 VSS.n11665 VSS.n11664 146.25
R4756 VSS.n11664 VSS.n11663 146.25
R4757 VSS.n11662 VSS.n11661 146.25
R4758 VSS.n11661 VSS.n11660 146.25
R4759 VSS.n11659 VSS.n11658 146.25
R4760 VSS.n11658 VSS.n11657 146.25
R4761 VSS.n11656 VSS.n11655 146.25
R4762 VSS.n11655 VSS.n11654 146.25
R4763 VSS.n11653 VSS.n11652 146.25
R4764 VSS.n11652 VSS.n11651 146.25
R4765 VSS.n11650 VSS.n11649 146.25
R4766 VSS.n11649 VSS.n11648 146.25
R4767 VSS.n11647 VSS.n11646 146.25
R4768 VSS.n11646 VSS.n11645 146.25
R4769 VSS.n11680 VSS.n11679 146.25
R4770 VSS.n11679 VSS.n11678 146.25
R4771 VSS.n11594 VSS.n11593 146.25
R4772 VSS.n11432 VSS.n11431 146.25
R4773 VSS.n11431 VSS.n11430 146.25
R4774 VSS.n11429 VSS.n11428 146.25
R4775 VSS.n11428 VSS.n11427 146.25
R4776 VSS.n11426 VSS.n11425 146.25
R4777 VSS.n11425 VSS.n11424 146.25
R4778 VSS.n11423 VSS.n11422 146.25
R4779 VSS.n11422 VSS.n11421 146.25
R4780 VSS.n11420 VSS.n11419 146.25
R4781 VSS.n11419 VSS.n11418 146.25
R4782 VSS.n11417 VSS.n11416 146.25
R4783 VSS.n11416 VSS.n11415 146.25
R4784 VSS.n11414 VSS.n11413 146.25
R4785 VSS.n11413 VSS.n11412 146.25
R4786 VSS.n11411 VSS.n11410 146.25
R4787 VSS.n11410 VSS.n11409 146.25
R4788 VSS.n11408 VSS.n11407 146.25
R4789 VSS.n11407 VSS.n11406 146.25
R4790 VSS.n11405 VSS.n11404 146.25
R4791 VSS.n11404 VSS.n11403 146.25
R4792 VSS.n11402 VSS.n11401 146.25
R4793 VSS.n11401 VSS.n11400 146.25
R4794 VSS.n11435 VSS.n11434 146.25
R4795 VSS.n11434 VSS.n11433 146.25
R4796 VSS.n11350 VSS.n11349 146.25
R4797 VSS.n11189 VSS.n11188 146.25
R4798 VSS.n11188 VSS.n11187 146.25
R4799 VSS.n11186 VSS.n11185 146.25
R4800 VSS.n11185 VSS.n11184 146.25
R4801 VSS.n11183 VSS.n11182 146.25
R4802 VSS.n11182 VSS.n11181 146.25
R4803 VSS.n11180 VSS.n11179 146.25
R4804 VSS.n11179 VSS.n11178 146.25
R4805 VSS.n11177 VSS.n11176 146.25
R4806 VSS.n11176 VSS.n11175 146.25
R4807 VSS.n11174 VSS.n11173 146.25
R4808 VSS.n11173 VSS.n11172 146.25
R4809 VSS.n11171 VSS.n11170 146.25
R4810 VSS.n11170 VSS.n11169 146.25
R4811 VSS.n11168 VSS.n11167 146.25
R4812 VSS.n11167 VSS.n11166 146.25
R4813 VSS.n11165 VSS.n11164 146.25
R4814 VSS.n11164 VSS.n11163 146.25
R4815 VSS.n11162 VSS.n11161 146.25
R4816 VSS.n11161 VSS.n11160 146.25
R4817 VSS.n11159 VSS.n11158 146.25
R4818 VSS.n11158 VSS.n11157 146.25
R4819 VSS.n11192 VSS.n11191 146.25
R4820 VSS.n11191 VSS.n11190 146.25
R4821 VSS.n11106 VSS.n11105 146.25
R4822 VSS.n10944 VSS.n10943 146.25
R4823 VSS.n10943 VSS.n10942 146.25
R4824 VSS.n10941 VSS.n10940 146.25
R4825 VSS.n10940 VSS.n10939 146.25
R4826 VSS.n10938 VSS.n10937 146.25
R4827 VSS.n10937 VSS.n10936 146.25
R4828 VSS.n10935 VSS.n10934 146.25
R4829 VSS.n10934 VSS.n10933 146.25
R4830 VSS.n10932 VSS.n10931 146.25
R4831 VSS.n10931 VSS.n10930 146.25
R4832 VSS.n10929 VSS.n10928 146.25
R4833 VSS.n10928 VSS.n10927 146.25
R4834 VSS.n10926 VSS.n10925 146.25
R4835 VSS.n10925 VSS.n10924 146.25
R4836 VSS.n10923 VSS.n10922 146.25
R4837 VSS.n10922 VSS.n10921 146.25
R4838 VSS.n10920 VSS.n10919 146.25
R4839 VSS.n10919 VSS.n10918 146.25
R4840 VSS.n10917 VSS.n10916 146.25
R4841 VSS.n10916 VSS.n10915 146.25
R4842 VSS.n10914 VSS.n10913 146.25
R4843 VSS.n10913 VSS.n10912 146.25
R4844 VSS.n10947 VSS.n10946 146.25
R4845 VSS.n10946 VSS.n10945 146.25
R4846 VSS.n10850 VSS.n10849 146.25
R4847 VSS.n8988 VSS.n8987 146.25
R4848 VSS.n8987 VSS.n8986 146.25
R4849 VSS.n8985 VSS.n8984 146.25
R4850 VSS.n8984 VSS.n8983 146.25
R4851 VSS.n8982 VSS.n8981 146.25
R4852 VSS.n8981 VSS.n8980 146.25
R4853 VSS.n8979 VSS.n8978 146.25
R4854 VSS.n8978 VSS.n8977 146.25
R4855 VSS.n8976 VSS.n8975 146.25
R4856 VSS.n8975 VSS.n8974 146.25
R4857 VSS.n8973 VSS.n8972 146.25
R4858 VSS.n8972 VSS.n8971 146.25
R4859 VSS.n8970 VSS.n8969 146.25
R4860 VSS.n8969 VSS.n8968 146.25
R4861 VSS.n8967 VSS.n8966 146.25
R4862 VSS.n8966 VSS.n8965 146.25
R4863 VSS.n8964 VSS.n8963 146.25
R4864 VSS.n8963 VSS.n8962 146.25
R4865 VSS.n8961 VSS.n8960 146.25
R4866 VSS.n8960 VSS.n8959 146.25
R4867 VSS.n8958 VSS.n8957 146.25
R4868 VSS.n8957 VSS.n8956 146.25
R4869 VSS.n8991 VSS.n8990 146.25
R4870 VSS.n8990 VSS.n8989 146.25
R4871 VSS.n8894 VSS.n8893 146.25
R4872 VSS.n8733 VSS.n8732 146.25
R4873 VSS.n8732 VSS.n8731 146.25
R4874 VSS.n8730 VSS.n8729 146.25
R4875 VSS.n8729 VSS.n8728 146.25
R4876 VSS.n8727 VSS.n8726 146.25
R4877 VSS.n8726 VSS.n8725 146.25
R4878 VSS.n8724 VSS.n8723 146.25
R4879 VSS.n8723 VSS.n8722 146.25
R4880 VSS.n8721 VSS.n8720 146.25
R4881 VSS.n8720 VSS.n8719 146.25
R4882 VSS.n8718 VSS.n8717 146.25
R4883 VSS.n8717 VSS.n8716 146.25
R4884 VSS.n8715 VSS.n8714 146.25
R4885 VSS.n8714 VSS.n8713 146.25
R4886 VSS.n8712 VSS.n8711 146.25
R4887 VSS.n8711 VSS.n8710 146.25
R4888 VSS.n8709 VSS.n8708 146.25
R4889 VSS.n8708 VSS.n8707 146.25
R4890 VSS.n8706 VSS.n8705 146.25
R4891 VSS.n8705 VSS.n8704 146.25
R4892 VSS.n8703 VSS.n8702 146.25
R4893 VSS.n8702 VSS.n8701 146.25
R4894 VSS.n8736 VSS.n8735 146.25
R4895 VSS.n8735 VSS.n8734 146.25
R4896 VSS.n8650 VSS.n8649 146.25
R4897 VSS.n8488 VSS.n8487 146.25
R4898 VSS.n8487 VSS.n8486 146.25
R4899 VSS.n8485 VSS.n8484 146.25
R4900 VSS.n8484 VSS.n8483 146.25
R4901 VSS.n8482 VSS.n8481 146.25
R4902 VSS.n8481 VSS.n8480 146.25
R4903 VSS.n8479 VSS.n8478 146.25
R4904 VSS.n8478 VSS.n8477 146.25
R4905 VSS.n8476 VSS.n8475 146.25
R4906 VSS.n8475 VSS.n8474 146.25
R4907 VSS.n8473 VSS.n8472 146.25
R4908 VSS.n8472 VSS.n8471 146.25
R4909 VSS.n8470 VSS.n8469 146.25
R4910 VSS.n8469 VSS.n8468 146.25
R4911 VSS.n8467 VSS.n8466 146.25
R4912 VSS.n8466 VSS.n8465 146.25
R4913 VSS.n8464 VSS.n8463 146.25
R4914 VSS.n8463 VSS.n8462 146.25
R4915 VSS.n8461 VSS.n8460 146.25
R4916 VSS.n8460 VSS.n8459 146.25
R4917 VSS.n8458 VSS.n8457 146.25
R4918 VSS.n8457 VSS.n8456 146.25
R4919 VSS.n8491 VSS.n8490 146.25
R4920 VSS.n8490 VSS.n8489 146.25
R4921 VSS.n8406 VSS.n8405 146.25
R4922 VSS.n8245 VSS.n8244 146.25
R4923 VSS.n8244 VSS.n8243 146.25
R4924 VSS.n8242 VSS.n8241 146.25
R4925 VSS.n8241 VSS.n8240 146.25
R4926 VSS.n8239 VSS.n8238 146.25
R4927 VSS.n8238 VSS.n8237 146.25
R4928 VSS.n8236 VSS.n8235 146.25
R4929 VSS.n8235 VSS.n8234 146.25
R4930 VSS.n8233 VSS.n8232 146.25
R4931 VSS.n8232 VSS.n8231 146.25
R4932 VSS.n8230 VSS.n8229 146.25
R4933 VSS.n8229 VSS.n8228 146.25
R4934 VSS.n8227 VSS.n8226 146.25
R4935 VSS.n8226 VSS.n8225 146.25
R4936 VSS.n8224 VSS.n8223 146.25
R4937 VSS.n8223 VSS.n8222 146.25
R4938 VSS.n8221 VSS.n8220 146.25
R4939 VSS.n8220 VSS.n8219 146.25
R4940 VSS.n8218 VSS.n8217 146.25
R4941 VSS.n8217 VSS.n8216 146.25
R4942 VSS.n8215 VSS.n8214 146.25
R4943 VSS.n8214 VSS.n8213 146.25
R4944 VSS.n8248 VSS.n8247 146.25
R4945 VSS.n8247 VSS.n8246 146.25
R4946 VSS.n8162 VSS.n8161 146.25
R4947 VSS.n8000 VSS.n7999 146.25
R4948 VSS.n7999 VSS.n7998 146.25
R4949 VSS.n7997 VSS.n7996 146.25
R4950 VSS.n7996 VSS.n7995 146.25
R4951 VSS.n7994 VSS.n7993 146.25
R4952 VSS.n7993 VSS.n7992 146.25
R4953 VSS.n7991 VSS.n7990 146.25
R4954 VSS.n7990 VSS.n7989 146.25
R4955 VSS.n7988 VSS.n7987 146.25
R4956 VSS.n7987 VSS.n7986 146.25
R4957 VSS.n7985 VSS.n7984 146.25
R4958 VSS.n7984 VSS.n7983 146.25
R4959 VSS.n7982 VSS.n7981 146.25
R4960 VSS.n7981 VSS.n7980 146.25
R4961 VSS.n7979 VSS.n7978 146.25
R4962 VSS.n7978 VSS.n7977 146.25
R4963 VSS.n7976 VSS.n7975 146.25
R4964 VSS.n7975 VSS.n7974 146.25
R4965 VSS.n7973 VSS.n7972 146.25
R4966 VSS.n7972 VSS.n7971 146.25
R4967 VSS.n7970 VSS.n7969 146.25
R4968 VSS.n7969 VSS.n7968 146.25
R4969 VSS.n8003 VSS.n8002 146.25
R4970 VSS.n8002 VSS.n8001 146.25
R4971 VSS.n7918 VSS.n7917 146.25
R4972 VSS.n7757 VSS.n7756 146.25
R4973 VSS.n7756 VSS.n7755 146.25
R4974 VSS.n7754 VSS.n7753 146.25
R4975 VSS.n7753 VSS.n7752 146.25
R4976 VSS.n7751 VSS.n7750 146.25
R4977 VSS.n7750 VSS.n7749 146.25
R4978 VSS.n7748 VSS.n7747 146.25
R4979 VSS.n7747 VSS.n7746 146.25
R4980 VSS.n7745 VSS.n7744 146.25
R4981 VSS.n7744 VSS.n7743 146.25
R4982 VSS.n7742 VSS.n7741 146.25
R4983 VSS.n7741 VSS.n7740 146.25
R4984 VSS.n7739 VSS.n7738 146.25
R4985 VSS.n7738 VSS.n7737 146.25
R4986 VSS.n7736 VSS.n7735 146.25
R4987 VSS.n7735 VSS.n7734 146.25
R4988 VSS.n7733 VSS.n7732 146.25
R4989 VSS.n7732 VSS.n7731 146.25
R4990 VSS.n7730 VSS.n7729 146.25
R4991 VSS.n7729 VSS.n7728 146.25
R4992 VSS.n7727 VSS.n7726 146.25
R4993 VSS.n7726 VSS.n7725 146.25
R4994 VSS.n7760 VSS.n7759 146.25
R4995 VSS.n7759 VSS.n7758 146.25
R4996 VSS.n7674 VSS.n7673 146.25
R4997 VSS.n7512 VSS.n7511 146.25
R4998 VSS.n7511 VSS.n7510 146.25
R4999 VSS.n7509 VSS.n7508 146.25
R5000 VSS.n7508 VSS.n7507 146.25
R5001 VSS.n7506 VSS.n7505 146.25
R5002 VSS.n7505 VSS.n7504 146.25
R5003 VSS.n7503 VSS.n7502 146.25
R5004 VSS.n7502 VSS.n7501 146.25
R5005 VSS.n7500 VSS.n7499 146.25
R5006 VSS.n7499 VSS.n7498 146.25
R5007 VSS.n7497 VSS.n7496 146.25
R5008 VSS.n7496 VSS.n7495 146.25
R5009 VSS.n7494 VSS.n7493 146.25
R5010 VSS.n7493 VSS.n7492 146.25
R5011 VSS.n7491 VSS.n7490 146.25
R5012 VSS.n7490 VSS.n7489 146.25
R5013 VSS.n7488 VSS.n7487 146.25
R5014 VSS.n7487 VSS.n7486 146.25
R5015 VSS.n7485 VSS.n7484 146.25
R5016 VSS.n7484 VSS.n7483 146.25
R5017 VSS.n7482 VSS.n7481 146.25
R5018 VSS.n7481 VSS.n7480 146.25
R5019 VSS.n7515 VSS.n7514 146.25
R5020 VSS.n7514 VSS.n7513 146.25
R5021 VSS.n7418 VSS.n7417 146.25
R5022 VSS.n1275 VSS.n1274 146.25
R5023 VSS.n1276 VSS.n1275 146.25
R5024 VSS.n647 VSS.n646 146.25
R5025 VSS.n1277 VSS.n647 146.25
R5026 VSS.n1280 VSS.n1279 146.25
R5027 VSS.n1279 VSS.n1278 146.25
R5028 VSS.n1281 VSS.n645 146.25
R5029 VSS.n645 VSS.n644 146.25
R5030 VSS.n1283 VSS.n1282 146.25
R5031 VSS.n1284 VSS.n1283 146.25
R5032 VSS.n643 VSS.n642 146.25
R5033 VSS.n1285 VSS.n643 146.25
R5034 VSS.n1288 VSS.n1287 146.25
R5035 VSS.n1287 VSS.n1286 146.25
R5036 VSS.n1289 VSS.n641 146.25
R5037 VSS.n641 VSS.n640 146.25
R5038 VSS.n1291 VSS.n1290 146.25
R5039 VSS.n1292 VSS.n1291 146.25
R5040 VSS.n639 VSS.n638 146.25
R5041 VSS.n1293 VSS.n639 146.25
R5042 VSS.n1296 VSS.n1295 146.25
R5043 VSS.n1295 VSS.n1294 146.25
R5044 VSS.n1273 VSS.n649 146.25
R5045 VSS.n649 VSS.n648 146.25
R5046 VSS.n1272 VSS.n1271 146.25
R5047 VSS.n1271 VSS.n1270 146.25
R5048 VSS.n912 VSS.n911 146.25
R5049 VSS.n911 VSS.n910 146.25
R5050 VSS.n887 VSS.n886 146.25
R5051 VSS.n909 VSS.n887 146.25
R5052 VSS.n907 VSS.n906 146.25
R5053 VSS.n908 VSS.n907 146.25
R5054 VSS.n905 VSS.n889 146.25
R5055 VSS.n889 VSS.n888 146.25
R5056 VSS.n904 VSS.n903 146.25
R5057 VSS.n903 VSS.n902 146.25
R5058 VSS.n891 VSS.n890 146.25
R5059 VSS.n901 VSS.n891 146.25
R5060 VSS.n899 VSS.n898 146.25
R5061 VSS.n900 VSS.n899 146.25
R5062 VSS.n897 VSS.n893 146.25
R5063 VSS.n893 VSS.n892 146.25
R5064 VSS.n896 VSS.n895 146.25
R5065 VSS.n895 VSS.n894 146.25
R5066 VSS.n623 VSS.n621 146.25
R5067 VSS.n621 VSS.n620 146.25
R5068 VSS.n1324 VSS.n1323 146.25
R5069 VSS.n1325 VSS.n1324 146.25
R5070 VSS.n913 VSS.n718 146.25
R5071 VSS.n718 VSS.n716 146.25
R5072 VSS.n915 VSS.n914 146.25
R5073 VSS.n916 VSS.n915 146.25
R5074 VSS.n5695 VSS.n5694 146.25
R5075 VSS.n5696 VSS.n5695 146.25
R5076 VSS.n5693 VSS.n596 146.25
R5077 VSS.n596 VSS.n595 146.25
R5078 VSS.n5692 VSS.n5691 146.25
R5079 VSS.n5691 VSS.n5690 146.25
R5080 VSS.n598 VSS.n597 146.25
R5081 VSS.n5689 VSS.n598 146.25
R5082 VSS.n5687 VSS.n5686 146.25
R5083 VSS.n5688 VSS.n5687 146.25
R5084 VSS.n5685 VSS.n600 146.25
R5085 VSS.n600 VSS.n599 146.25
R5086 VSS.n5684 VSS.n5683 146.25
R5087 VSS.n5683 VSS.n5682 146.25
R5088 VSS.n602 VSS.n601 146.25
R5089 VSS.n5681 VSS.n602 146.25
R5090 VSS.n5679 VSS.n5678 146.25
R5091 VSS.n5680 VSS.n5679 146.25
R5092 VSS.n5677 VSS.n604 146.25
R5093 VSS.n604 VSS.n603 146.25
R5094 VSS.n5676 VSS.n5675 146.25
R5095 VSS.n5675 VSS.n5674 146.25
R5096 VSS.n593 VSS.n591 146.25
R5097 VSS.n5697 VSS.n593 146.25
R5098 VSS.n5700 VSS.n5699 146.25
R5099 VSS.n5699 VSS.n5698 146.25
R5100 VSS.n1377 VSS.n1376 146.25
R5101 VSS.n5622 VSS.n1377 146.25
R5102 VSS.n5625 VSS.n5624 146.25
R5103 VSS.n5624 VSS.n5623 146.25
R5104 VSS.n5626 VSS.n1375 146.25
R5105 VSS.n1375 VSS.n1374 146.25
R5106 VSS.n5628 VSS.n5627 146.25
R5107 VSS.n5629 VSS.n5628 146.25
R5108 VSS.n1373 VSS.n1372 146.25
R5109 VSS.n5630 VSS.n1373 146.25
R5110 VSS.n5633 VSS.n5632 146.25
R5111 VSS.n5632 VSS.n5631 146.25
R5112 VSS.n5634 VSS.n1371 146.25
R5113 VSS.n1371 VSS.n1370 146.25
R5114 VSS.n5637 VSS.n5636 146.25
R5115 VSS.n5638 VSS.n5637 146.25
R5116 VSS.n5635 VSS.n1369 146.25
R5117 VSS.n5639 VSS.n1369 146.25
R5118 VSS.n5641 VSS.n1368 146.25
R5119 VSS.n5641 VSS.n5640 146.25
R5120 VSS.n5643 VSS.n5642 146.25
R5121 VSS.n5642 VSS.n1363 146.25
R5122 VSS.n5620 VSS.n5619 146.25
R5123 VSS.n5621 VSS.n5620 146.25
R5124 VSS.n5618 VSS.n1379 146.25
R5125 VSS.n1379 VSS.n1378 146.25
R5126 VSS.n5487 VSS.n5486 146.25
R5127 VSS.n5488 VSS.n5487 146.25
R5128 VSS.n5485 VSS.n1451 146.25
R5129 VSS.n1451 VSS.n1450 146.25
R5130 VSS.n5484 VSS.n5483 146.25
R5131 VSS.n5483 VSS.n5482 146.25
R5132 VSS.n1453 VSS.n1452 146.25
R5133 VSS.n5481 VSS.n1453 146.25
R5134 VSS.n5479 VSS.n5478 146.25
R5135 VSS.n5480 VSS.n5479 146.25
R5136 VSS.n5477 VSS.n1455 146.25
R5137 VSS.n1455 VSS.n1454 146.25
R5138 VSS.n5476 VSS.n5475 146.25
R5139 VSS.n5475 VSS.n5474 146.25
R5140 VSS.n1457 VSS.n1456 146.25
R5141 VSS.n5473 VSS.n1457 146.25
R5142 VSS.n5471 VSS.n5470 146.25
R5143 VSS.n5472 VSS.n5471 146.25
R5144 VSS.n5469 VSS.n1459 146.25
R5145 VSS.n1459 VSS.n1458 146.25
R5146 VSS.n5468 VSS.n5467 146.25
R5147 VSS.n5467 VSS.n5466 146.25
R5148 VSS.n1449 VSS.n1448 146.25
R5149 VSS.n5489 VSS.n1449 146.25
R5150 VSS.n5492 VSS.n5491 146.25
R5151 VSS.n5491 VSS.n5490 146.25
R5152 VSS.n1518 VSS.n1517 146.25
R5153 VSS.n5414 VSS.n1518 146.25
R5154 VSS.n5417 VSS.n5416 146.25
R5155 VSS.n5416 VSS.n5415 146.25
R5156 VSS.n5418 VSS.n1516 146.25
R5157 VSS.n1516 VSS.n1515 146.25
R5158 VSS.n5420 VSS.n5419 146.25
R5159 VSS.n5421 VSS.n5420 146.25
R5160 VSS.n1514 VSS.n1513 146.25
R5161 VSS.n5422 VSS.n1514 146.25
R5162 VSS.n5425 VSS.n5424 146.25
R5163 VSS.n5424 VSS.n5423 146.25
R5164 VSS.n5426 VSS.n1512 146.25
R5165 VSS.n1512 VSS.n1511 146.25
R5166 VSS.n5429 VSS.n5428 146.25
R5167 VSS.n5430 VSS.n5429 146.25
R5168 VSS.n5427 VSS.n1510 146.25
R5169 VSS.n5431 VSS.n1510 146.25
R5170 VSS.n5433 VSS.n1509 146.25
R5171 VSS.n5433 VSS.n5432 146.25
R5172 VSS.n5435 VSS.n5434 146.25
R5173 VSS.n5434 VSS.n1504 146.25
R5174 VSS.n5412 VSS.n5411 146.25
R5175 VSS.n5413 VSS.n5412 146.25
R5176 VSS.n5410 VSS.n1520 146.25
R5177 VSS.n1520 VSS.n1519 146.25
R5178 VSS.n4754 VSS.n4753 146.25
R5179 VSS.n4755 VSS.n4754 146.25
R5180 VSS.n4752 VSS.n4730 146.25
R5181 VSS.n4730 VSS.n4729 146.25
R5182 VSS.n4751 VSS.n4750 146.25
R5183 VSS.n4750 VSS.n4749 146.25
R5184 VSS.n4732 VSS.n4731 146.25
R5185 VSS.n4748 VSS.n4732 146.25
R5186 VSS.n4746 VSS.n4745 146.25
R5187 VSS.n4747 VSS.n4746 146.25
R5188 VSS.n4744 VSS.n4734 146.25
R5189 VSS.n4734 VSS.n4733 146.25
R5190 VSS.n4743 VSS.n4742 146.25
R5191 VSS.n4742 VSS.n4741 146.25
R5192 VSS.n4736 VSS.n4735 146.25
R5193 VSS.n4740 VSS.n4736 146.25
R5194 VSS.n4738 VSS.n4737 146.25
R5195 VSS.n4739 VSS.n4738 146.25
R5196 VSS.n3125 VSS.n3124 146.25
R5197 VSS.n3127 VSS.n3125 146.25
R5198 VSS.n5079 VSS.n5078 146.25
R5199 VSS.n5078 VSS.n5077 146.25
R5200 VSS.n4728 VSS.n4727 146.25
R5201 VSS.n4756 VSS.n4728 146.25
R5202 VSS.n4759 VSS.n4758 146.25
R5203 VSS.n4758 VSS.n4757 146.25
R5204 VSS.n5029 VSS.n5028 146.25
R5205 VSS.n5028 VSS.n5027 146.25
R5206 VSS.n5030 VSS.n3150 146.25
R5207 VSS.n3150 VSS.n3149 146.25
R5208 VSS.n5032 VSS.n5031 146.25
R5209 VSS.n5033 VSS.n5032 146.25
R5210 VSS.n3148 VSS.n3147 146.25
R5211 VSS.n5034 VSS.n3148 146.25
R5212 VSS.n5037 VSS.n5036 146.25
R5213 VSS.n5036 VSS.n5035 146.25
R5214 VSS.n5038 VSS.n3146 146.25
R5215 VSS.n3146 VSS.n3145 146.25
R5216 VSS.n5040 VSS.n5039 146.25
R5217 VSS.n5041 VSS.n5040 146.25
R5218 VSS.n3144 VSS.n3143 146.25
R5219 VSS.n5042 VSS.n3144 146.25
R5220 VSS.n5045 VSS.n5044 146.25
R5221 VSS.n5044 VSS.n5043 146.25
R5222 VSS.n5046 VSS.n3142 146.25
R5223 VSS.n3142 VSS.n3141 146.25
R5224 VSS.n5048 VSS.n5047 146.25
R5225 VSS.n5049 VSS.n5048 146.25
R5226 VSS.n3152 VSS.n3151 146.25
R5227 VSS.n5026 VSS.n3152 146.25
R5228 VSS.n5024 VSS.n5023 146.25
R5229 VSS.n5025 VSS.n5024 146.25
R5230 VSS.n4525 VSS.n4524 146.25
R5231 VSS.n4526 VSS.n4525 146.25
R5232 VSS.n4523 VSS.n3231 146.25
R5233 VSS.n3231 VSS.n3230 146.25
R5234 VSS.n4522 VSS.n4521 146.25
R5235 VSS.n4521 VSS.n4520 146.25
R5236 VSS.n3234 VSS.n3233 146.25
R5237 VSS.n4519 VSS.n3234 146.25
R5238 VSS.n4517 VSS.n4516 146.25
R5239 VSS.n4518 VSS.n4517 146.25
R5240 VSS.n4515 VSS.n3236 146.25
R5241 VSS.n3236 VSS.n3235 146.25
R5242 VSS.n4514 VSS.n4513 146.25
R5243 VSS.n4513 VSS.n4512 146.25
R5244 VSS.n3238 VSS.n3237 146.25
R5245 VSS.n4511 VSS.n3238 146.25
R5246 VSS.n4509 VSS.n4508 146.25
R5247 VSS.n4510 VSS.n4509 146.25
R5248 VSS.n4507 VSS.n3240 146.25
R5249 VSS.n3240 VSS.n3239 146.25
R5250 VSS.n4506 VSS.n4505 146.25
R5251 VSS.n4505 VSS.n4504 146.25
R5252 VSS.n3232 VSS.n3229 146.25
R5253 VSS.n4527 VSS.n3229 146.25
R5254 VSS.n4529 VSS.n3220 146.25
R5255 VSS.n4529 VSS.n4528 146.25
R5256 VSS.n4164 VSS.n4163 146.25
R5257 VSS.n4165 VSS.n4164 146.25
R5258 VSS.n4162 VSS.n4140 146.25
R5259 VSS.n4140 VSS.n4139 146.25
R5260 VSS.n4161 VSS.n4160 146.25
R5261 VSS.n4160 VSS.n4159 146.25
R5262 VSS.n4142 VSS.n4141 146.25
R5263 VSS.n4158 VSS.n4142 146.25
R5264 VSS.n4156 VSS.n4155 146.25
R5265 VSS.n4157 VSS.n4156 146.25
R5266 VSS.n4154 VSS.n4144 146.25
R5267 VSS.n4144 VSS.n4143 146.25
R5268 VSS.n4153 VSS.n4152 146.25
R5269 VSS.n4152 VSS.n4151 146.25
R5270 VSS.n4146 VSS.n4145 146.25
R5271 VSS.n4150 VSS.n4146 146.25
R5272 VSS.n4148 VSS.n4147 146.25
R5273 VSS.n4149 VSS.n4148 146.25
R5274 VSS.n3294 VSS.n3292 146.25
R5275 VSS.n3292 VSS.n3291 146.25
R5276 VSS.n4476 VSS.n4475 146.25
R5277 VSS.n4477 VSS.n4476 146.25
R5278 VSS.n4138 VSS.n4137 146.25
R5279 VSS.n4166 VSS.n4138 146.25
R5280 VSS.n4169 VSS.n4168 146.25
R5281 VSS.n4168 VSS.n4167 146.25
R5282 VSS.n4426 VSS.n4425 146.25
R5283 VSS.n4427 VSS.n4426 146.25
R5284 VSS.n3317 VSS.n3316 146.25
R5285 VSS.n4428 VSS.n3317 146.25
R5286 VSS.n4431 VSS.n4430 146.25
R5287 VSS.n4430 VSS.n4429 146.25
R5288 VSS.n4432 VSS.n3315 146.25
R5289 VSS.n3315 VSS.n3314 146.25
R5290 VSS.n4434 VSS.n4433 146.25
R5291 VSS.n4435 VSS.n4434 146.25
R5292 VSS.n3313 VSS.n3312 146.25
R5293 VSS.n4436 VSS.n3313 146.25
R5294 VSS.n4439 VSS.n4438 146.25
R5295 VSS.n4438 VSS.n4437 146.25
R5296 VSS.n4440 VSS.n3311 146.25
R5297 VSS.n3311 VSS.n3310 146.25
R5298 VSS.n4442 VSS.n4441 146.25
R5299 VSS.n4443 VSS.n4442 146.25
R5300 VSS.n3309 VSS.n3308 146.25
R5301 VSS.n4444 VSS.n3309 146.25
R5302 VSS.n4447 VSS.n4446 146.25
R5303 VSS.n4446 VSS.n4445 146.25
R5304 VSS.n4424 VSS.n3319 146.25
R5305 VSS.n3319 VSS.n3318 146.25
R5306 VSS.n4423 VSS.n4422 146.25
R5307 VSS.n4422 VSS.n4421 146.25
R5308 VSS.n3396 VSS.n3393 146.25
R5309 VSS.n3946 VSS.n3393 146.25
R5310 VSS.n3944 VSS.n3943 146.25
R5311 VSS.n3945 VSS.n3944 146.25
R5312 VSS.n3942 VSS.n3395 146.25
R5313 VSS.n3395 VSS.n3394 146.25
R5314 VSS.n3941 VSS.n3940 146.25
R5315 VSS.n3940 VSS.n3939 146.25
R5316 VSS.n3398 VSS.n3397 146.25
R5317 VSS.n3938 VSS.n3398 146.25
R5318 VSS.n3936 VSS.n3935 146.25
R5319 VSS.n3937 VSS.n3936 146.25
R5320 VSS.n3934 VSS.n3400 146.25
R5321 VSS.n3400 VSS.n3399 146.25
R5322 VSS.n3933 VSS.n3932 146.25
R5323 VSS.n3932 VSS.n3931 146.25
R5324 VSS.n3402 VSS.n3401 146.25
R5325 VSS.n3930 VSS.n3402 146.25
R5326 VSS.n3928 VSS.n3927 146.25
R5327 VSS.n3929 VSS.n3928 146.25
R5328 VSS.n3926 VSS.n3404 146.25
R5329 VSS.n3404 VSS.n3403 146.25
R5330 VSS.n3948 VSS.n3392 146.25
R5331 VSS.n3948 VSS.n3947 146.25
R5332 VSS.n3950 VSS.n3949 146.25
R5333 VSS.n3949 VSS.n3385 146.25
R5334 VSS.n3552 VSS.n3551 146.25
R5335 VSS.n3553 VSS.n3552 146.25
R5336 VSS.n3550 VSS.n3528 146.25
R5337 VSS.n3528 VSS.n3527 146.25
R5338 VSS.n3549 VSS.n3548 146.25
R5339 VSS.n3548 VSS.n3547 146.25
R5340 VSS.n3530 VSS.n3529 146.25
R5341 VSS.n3546 VSS.n3530 146.25
R5342 VSS.n3544 VSS.n3543 146.25
R5343 VSS.n3545 VSS.n3544 146.25
R5344 VSS.n3542 VSS.n3532 146.25
R5345 VSS.n3532 VSS.n3531 146.25
R5346 VSS.n3541 VSS.n3540 146.25
R5347 VSS.n3540 VSS.n3539 146.25
R5348 VSS.n3534 VSS.n3533 146.25
R5349 VSS.n3538 VSS.n3534 146.25
R5350 VSS.n3536 VSS.n3535 146.25
R5351 VSS.n3537 VSS.n3536 146.25
R5352 VSS.n3421 VSS.n3420 146.25
R5353 VSS.n3423 VSS.n3421 146.25
R5354 VSS.n3864 VSS.n3863 146.25
R5355 VSS.n3863 VSS.n3862 146.25
R5356 VSS.n3526 VSS.n3525 146.25
R5357 VSS.n3554 VSS.n3526 146.25
R5358 VSS.n3557 VSS.n3556 146.25
R5359 VSS.n3556 VSS.n3555 146.25
R5360 VSS.n14729 VSS.n14725 142.386
R5361 VSS.n14742 VSS.n14741 142.386
R5362 VSS.n15229 VSS.n15225 142.386
R5363 VSS.n15242 VSS.n15241 142.386
R5364 VSS.n14985 VSS.n14981 142.386
R5365 VSS.n14998 VSS.n14997 142.386
R5366 VSS.n15717 VSS.n15713 142.386
R5367 VSS.n15730 VSS.n15729 142.386
R5368 VSS.n15473 VSS.n15469 142.386
R5369 VSS.n15486 VSS.n15485 142.386
R5370 VSS.n16205 VSS.n16201 142.386
R5371 VSS.n16218 VSS.n16217 142.386
R5372 VSS.n15961 VSS.n15957 142.386
R5373 VSS.n15974 VSS.n15973 142.386
R5374 VSS.n16461 VSS.n16457 142.386
R5375 VSS.n16474 VSS.n16473 142.386
R5376 VSS.n10778 VSS.n10774 142.386
R5377 VSS.n10791 VSS.n10790 142.386
R5378 VSS.n11278 VSS.n11274 142.386
R5379 VSS.n11291 VSS.n11290 142.386
R5380 VSS.n11034 VSS.n11030 142.386
R5381 VSS.n11047 VSS.n11046 142.386
R5382 VSS.n11766 VSS.n11762 142.386
R5383 VSS.n11779 VSS.n11778 142.386
R5384 VSS.n11522 VSS.n11518 142.386
R5385 VSS.n11535 VSS.n11534 142.386
R5386 VSS.n12254 VSS.n12250 142.386
R5387 VSS.n12267 VSS.n12266 142.386
R5388 VSS.n12010 VSS.n12006 142.386
R5389 VSS.n12023 VSS.n12022 142.386
R5390 VSS.n12510 VSS.n12506 142.386
R5391 VSS.n12523 VSS.n12522 142.386
R5392 VSS.n7346 VSS.n7342 142.386
R5393 VSS.n7359 VSS.n7358 142.386
R5394 VSS.n7846 VSS.n7842 142.386
R5395 VSS.n7859 VSS.n7858 142.386
R5396 VSS.n7602 VSS.n7598 142.386
R5397 VSS.n7615 VSS.n7614 142.386
R5398 VSS.n8334 VSS.n8330 142.386
R5399 VSS.n8347 VSS.n8346 142.386
R5400 VSS.n8090 VSS.n8086 142.386
R5401 VSS.n8103 VSS.n8102 142.386
R5402 VSS.n8822 VSS.n8818 142.386
R5403 VSS.n8835 VSS.n8834 142.386
R5404 VSS.n8578 VSS.n8574 142.386
R5405 VSS.n8591 VSS.n8590 142.386
R5406 VSS.n9078 VSS.n9074 142.386
R5407 VSS.n9091 VSS.n9090 142.386
R5408 VSS.n5140 VSS.n1579 142.386
R5409 VSS.n5152 VSS.n1577 142.386
R5410 VSS.n5159 VSS.n1569 142.386
R5411 VSS.n5171 VSS.n1565 142.386
R5412 VSS.n5175 VSS.n1558 142.386
R5413 VSS.n5187 VSS.n1556 142.386
R5414 VSS.n5194 VSS.n1548 142.386
R5415 VSS.n5206 VSS.n1544 142.386
R5416 VSS.n5210 VSS.n1537 142.386
R5417 VSS.n5223 VSS.n1534 142.386
R5418 VSS.n5232 VSS.n1529 142.386
R5419 VSS.n5499 VSS.n1438 142.386
R5420 VSS.n5511 VSS.n1436 142.386
R5421 VSS.n5518 VSS.n1428 142.386
R5422 VSS.n5530 VSS.n1424 142.386
R5423 VSS.n5534 VSS.n1417 142.386
R5424 VSS.n5546 VSS.n1415 142.386
R5425 VSS.n5553 VSS.n1407 142.386
R5426 VSS.n5565 VSS.n1403 142.386
R5427 VSS.n5569 VSS.n1396 142.386
R5428 VSS.n5582 VSS.n1393 142.386
R5429 VSS.n5591 VSS.n1388 142.386
R5430 VSS.n5390 VSS.n5236 142.386
R5431 VSS.n5386 VSS.n5243 142.386
R5432 VSS.n5379 VSS.n5250 142.386
R5433 VSS.n5367 VSS.n5253 142.386
R5434 VSS.n5363 VSS.n5262 142.386
R5435 VSS.n5356 VSS.n5269 142.386
R5436 VSS.n5344 VSS.n5272 142.386
R5437 VSS.n5340 VSS.n5281 142.386
R5438 VSS.n5333 VSS.n5288 142.386
R5439 VSS.n5321 VSS.n5291 142.386
R5440 VSS.n5317 VSS.n5300 142.386
R5441 VSS.n785 VSS.n775 142.386
R5442 VSS.n797 VSS.n773 142.386
R5443 VSS.n804 VSS.n765 142.386
R5444 VSS.n816 VSS.n761 142.386
R5445 VSS.n820 VSS.n754 142.386
R5446 VSS.n832 VSS.n752 142.386
R5447 VSS.n839 VSS.n744 142.386
R5448 VSS.n851 VSS.n740 142.386
R5449 VSS.n855 VSS.n733 142.386
R5450 VSS.n867 VSS.n731 142.386
R5451 VSS.n874 VSS.n722 142.386
R5452 VSS.n5598 VSS.n5595 142.386
R5453 VSS.n5781 VSS.n524 142.386
R5454 VSS.n5769 VSS.n527 142.386
R5455 VSS.n5765 VSS.n536 142.386
R5456 VSS.n5758 VSS.n543 142.386
R5457 VSS.n5746 VSS.n546 142.386
R5458 VSS.n5742 VSS.n555 142.386
R5459 VSS.n5735 VSS.n562 142.386
R5460 VSS.n5723 VSS.n565 142.386
R5461 VSS.n5719 VSS.n574 142.386
R5462 VSS.n5712 VSS.n581 142.386
R5463 VSS.n928 VSS.n710 142.386
R5464 VSS.n932 VSS.n703 142.386
R5465 VSS.n944 VSS.n701 142.386
R5466 VSS.n951 VSS.n693 142.386
R5467 VSS.n963 VSS.n689 142.386
R5468 VSS.n967 VSS.n682 142.386
R5469 VSS.n979 VSS.n680 142.386
R5470 VSS.n986 VSS.n672 142.386
R5471 VSS.n998 VSS.n668 142.386
R5472 VSS.n1002 VSS.n661 142.386
R5473 VSS.n1014 VSS.n659 142.386
R5474 VSS.n1258 VSS.n1024 142.386
R5475 VSS.n1246 VSS.n1027 142.386
R5476 VSS.n1242 VSS.n1036 142.386
R5477 VSS.n1235 VSS.n1043 142.386
R5478 VSS.n1223 VSS.n1046 142.386
R5479 VSS.n1219 VSS.n1055 142.386
R5480 VSS.n1212 VSS.n1062 142.386
R5481 VSS.n1200 VSS.n1065 142.386
R5482 VSS.n1196 VSS.n1074 142.386
R5483 VSS.n1189 VSS.n1081 142.386
R5484 VSS.n1177 VSS.n1084 142.386
R5485 VSS.n3805 VSS.n3454 142.386
R5486 VSS.n3793 VSS.n3456 142.386
R5487 VSS.n3789 VSS.n3466 142.386
R5488 VSS.n3782 VSS.n3473 142.386
R5489 VSS.n3770 VSS.n3476 142.386
R5490 VSS.n3766 VSS.n3485 142.386
R5491 VSS.n3759 VSS.n3492 142.386
R5492 VSS.n3747 VSS.n3495 142.386
R5493 VSS.n3743 VSS.n3504 142.386
R5494 VSS.n3736 VSS.n3511 142.386
R5495 VSS.n3724 VSS.n3514 142.386
R5496 VSS.n3970 VSS.n3380 142.386
R5497 VSS.n3974 VSS.n3373 142.386
R5498 VSS.n3986 VSS.n3371 142.386
R5499 VSS.n3993 VSS.n3363 142.386
R5500 VSS.n4005 VSS.n3359 142.386
R5501 VSS.n4009 VSS.n3352 142.386
R5502 VSS.n4021 VSS.n3350 142.386
R5503 VSS.n4028 VSS.n3342 142.386
R5504 VSS.n4040 VSS.n3338 142.386
R5505 VSS.n4044 VSS.n3331 142.386
R5506 VSS.n4056 VSS.n3329 142.386
R5507 VSS.n3712 VSS.n3563 142.386
R5508 VSS.n3700 VSS.n3569 142.386
R5509 VSS.n3696 VSS.n3578 142.386
R5510 VSS.n3689 VSS.n3585 142.386
R5511 VSS.n3677 VSS.n3588 142.386
R5512 VSS.n3673 VSS.n3597 142.386
R5513 VSS.n3666 VSS.n3604 142.386
R5514 VSS.n3654 VSS.n3607 142.386
R5515 VSS.n3650 VSS.n3616 142.386
R5516 VSS.n3643 VSS.n3623 142.386
R5517 VSS.n3629 VSS.n3626 142.386
R5518 VSS.n4316 VSS.n4175 142.386
R5519 VSS.n4304 VSS.n4181 142.386
R5520 VSS.n4300 VSS.n4190 142.386
R5521 VSS.n4293 VSS.n4197 142.386
R5522 VSS.n4281 VSS.n4200 142.386
R5523 VSS.n4277 VSS.n4209 142.386
R5524 VSS.n4270 VSS.n4216 142.386
R5525 VSS.n4258 VSS.n4219 142.386
R5526 VSS.n4254 VSS.n4228 142.386
R5527 VSS.n4247 VSS.n4235 142.386
R5528 VSS.n4535 VSS.n3225 142.386
R5529 VSS.n4409 VSS.n4066 142.386
R5530 VSS.n4397 VSS.n4069 142.386
R5531 VSS.n4393 VSS.n4078 142.386
R5532 VSS.n4386 VSS.n4085 142.386
R5533 VSS.n4374 VSS.n4088 142.386
R5534 VSS.n4370 VSS.n4097 142.386
R5535 VSS.n4363 VSS.n4104 142.386
R5536 VSS.n4351 VSS.n4107 142.386
R5537 VSS.n4347 VSS.n4116 142.386
R5538 VSS.n4340 VSS.n4123 142.386
R5539 VSS.n4328 VSS.n4126 142.386
R5540 VSS.n5018 VSS.n4654 142.386
R5541 VSS.n5006 VSS.n4659 142.386
R5542 VSS.n5002 VSS.n4668 142.386
R5543 VSS.n4995 VSS.n4675 142.386
R5544 VSS.n4983 VSS.n4678 142.386
R5545 VSS.n4979 VSS.n4687 142.386
R5546 VSS.n4972 VSS.n4694 142.386
R5547 VSS.n4960 VSS.n4697 142.386
R5548 VSS.n4956 VSS.n4706 142.386
R5549 VSS.n4949 VSS.n4713 142.386
R5550 VSS.n4937 VSS.n4716 142.386
R5551 VSS.n4552 VSS.n3215 142.386
R5552 VSS.n4559 VSS.n3207 142.386
R5553 VSS.n4571 VSS.n3203 142.386
R5554 VSS.n4575 VSS.n3196 142.386
R5555 VSS.n4587 VSS.n3194 142.386
R5556 VSS.n4594 VSS.n3186 142.386
R5557 VSS.n4606 VSS.n3182 142.386
R5558 VSS.n4610 VSS.n3175 142.386
R5559 VSS.n4622 VSS.n3173 142.386
R5560 VSS.n4629 VSS.n3165 142.386
R5561 VSS.n4641 VSS.n3161 142.386
R5562 VSS.n4925 VSS.n4765 142.386
R5563 VSS.n4913 VSS.n4771 142.386
R5564 VSS.n4909 VSS.n4780 142.386
R5565 VSS.n4902 VSS.n4787 142.386
R5566 VSS.n4890 VSS.n4790 142.386
R5567 VSS.n4886 VSS.n4799 142.386
R5568 VSS.n4879 VSS.n4806 142.386
R5569 VSS.n4867 VSS.n4809 142.386
R5570 VSS.n4863 VSS.n4818 142.386
R5571 VSS.n4856 VSS.n4825 142.386
R5572 VSS.n4844 VSS.n4828 142.386
R5573 VSS.n379 VSS.n378 141.612
R5574 VSS.n436 VSS.n344 141.612
R5575 VSS.n18171 VSS.n18170 141.612
R5576 VSS.n18224 VSS.n18135 141.612
R5577 VSS.n375 VSS 130.062
R5578 VSS.n1164 VSS.n1093 126.781
R5579 VSS.n5127 VSS.n3098 126.781
R5580 VSS.n17879 VSS.n17792 126.781
R5581 VSS.n1651 VSS.n1586 124.831
R5582 VSS.n3813 VSS.n3447 124.831
R5583 VSS.n17851 VSS.n17806 124.831
R5584 VSS.n386 VSS.n385 109.655
R5585 VSS.n396 VSS.n392 109.655
R5586 VSS.n394 VSS.n362 109.655
R5587 VSS.n407 VSS.n405 109.655
R5588 VSS.n407 VSS.n406 109.655
R5589 VSS.n413 VSS.n412 109.655
R5590 VSS.n420 VSS.n419 109.655
R5591 VSS.n428 VSS.n426 109.655
R5592 VSS.n18178 VSS.n18177 109.655
R5593 VSS.n18188 VSS.n18184 109.655
R5594 VSS.n18186 VSS.n18154 109.655
R5595 VSS.n18199 VSS.n18197 109.655
R5596 VSS.n18199 VSS.n18198 109.655
R5597 VSS.n18205 VSS.n18204 109.655
R5598 VSS.n18213 VSS.n18212 109.655
R5599 VSS.n18222 VSS.n18139 109.655
R5600 VSS.n1507 VSS.n1503 97.524
R5601 VSS.n1366 VSS.n1362 97.524
R5602 VSS.n1490 VSS.n1461 97.524
R5603 VSS.n1320 VSS.n622 97.524
R5604 VSS.n1349 VSS.n606 97.524
R5605 VSS.n1118 VSS.n636 97.524
R5606 VSS.n3422 VSS.n3418 97.524
R5607 VSS.n4450 VSS.n3306 97.524
R5608 VSS.n3919 VSS.n3408 97.524
R5609 VSS.n3276 VSS.n3242 97.524
R5610 VSS.n3293 VSS.n3289 97.524
R5611 VSS.n5052 VSS.n3139 97.524
R5612 VSS.n3126 VSS.n3122 97.524
R5613 VSS.n18025 VSS 94.85
R5614 VSS.n2406 VSS.n2307 92.501
R5615 VSS.n2496 VSS.n2217 92.501
R5616 VSS.n2586 VSS.n2127 92.501
R5617 VSS.n2676 VSS.n2037 92.501
R5618 VSS.n2766 VSS.n1947 92.501
R5619 VSS.n2856 VSS.n1857 92.501
R5620 VSS.n2946 VSS.n1767 92.501
R5621 VSS.n3036 VSS.n1677 92.501
R5622 VSS.n6851 VSS.n6421 92.501
R5623 VSS.n6761 VSS.n6511 92.501
R5624 VSS.n6671 VSS.n6601 92.501
R5625 VSS.n14477 VSS.n14476 92.5
R5626 VSS.n14442 VSS.n14441 92.5
R5627 VSS.n14436 VSS.n14435 92.5
R5628 VSS.n14438 VSS.n14437 92.5
R5629 VSS.n14431 VSS.n14430 92.5
R5630 VSS.n14433 VSS.n14432 92.5
R5631 VSS.n14427 VSS.n14426 92.5
R5632 VSS.t10 VSS.n14440 92.5
R5633 VSS.n14310 VSS.n14309 92.5
R5634 VSS.n14297 VSS.n14296 92.5
R5635 VSS.n14262 VSS.n14261 92.5
R5636 VSS.n14256 VSS.n14255 92.5
R5637 VSS.n14258 VSS.n14257 92.5
R5638 VSS.n14251 VSS.n14250 92.5
R5639 VSS.n14253 VSS.n14252 92.5
R5640 VSS.n14247 VSS.n14246 92.5
R5641 VSS.t8 VSS.n14260 92.5
R5642 VSS.n14131 VSS.n14130 92.5
R5643 VSS.n17552 VSS.n17551 92.5
R5644 VSS.n17544 VSS.n17543 92.5
R5645 VSS.n17546 VSS.n17545 92.5
R5646 VSS.n17539 VSS.n17538 92.5
R5647 VSS.n17541 VSS.n17540 92.5
R5648 VSS.n17535 VSS.n17534 92.5
R5649 VSS.t6 VSS.n17533 92.5
R5650 VSS.n17384 VSS.n17383 92.5
R5651 VSS.n17376 VSS.n17375 92.5
R5652 VSS.n17378 VSS.n17377 92.5
R5653 VSS.n17371 VSS.n17370 92.5
R5654 VSS.n17373 VSS.n17372 92.5
R5655 VSS.n17367 VSS.n17366 92.5
R5656 VSS.t2 VSS.n17365 92.5
R5657 VSS.n17216 VSS.n17215 92.5
R5658 VSS.n17208 VSS.n17207 92.5
R5659 VSS.n17210 VSS.n17209 92.5
R5660 VSS.n17203 VSS.n17202 92.5
R5661 VSS.n17205 VSS.n17204 92.5
R5662 VSS.n17199 VSS.n17198 92.5
R5663 VSS.t4 VSS.n17197 92.5
R5664 VSS.n17048 VSS.n17047 92.5
R5665 VSS.n17040 VSS.n17039 92.5
R5666 VSS.n17042 VSS.n17041 92.5
R5667 VSS.n17035 VSS.n17034 92.5
R5668 VSS.n17037 VSS.n17036 92.5
R5669 VSS.n17031 VSS.n17030 92.5
R5670 VSS.t12 VSS.n17029 92.5
R5671 VSS.n16880 VSS.n16879 92.5
R5672 VSS.n16872 VSS.n16871 92.5
R5673 VSS.n16874 VSS.n16873 92.5
R5674 VSS.n16867 VSS.n16866 92.5
R5675 VSS.n16869 VSS.n16868 92.5
R5676 VSS.n16863 VSS.n16862 92.5
R5677 VSS.t14 VSS.n16861 92.5
R5678 VSS.n16712 VSS.n16711 92.5
R5679 VSS.n16704 VSS.n16703 92.5
R5680 VSS.n16706 VSS.n16705 92.5
R5681 VSS.n16699 VSS.n16698 92.5
R5682 VSS.n16701 VSS.n16700 92.5
R5683 VSS.n16695 VSS.n16694 92.5
R5684 VSS.t0 VSS.n16693 92.5
R5685 VSS.n14075 VSS.n14074 92.5
R5686 VSS.n14039 VSS.n14038 92.5
R5687 VSS.n14033 VSS.n14032 92.5
R5688 VSS.n14035 VSS.n14034 92.5
R5689 VSS.n14028 VSS.n14027 92.5
R5690 VSS.n14030 VSS.n14029 92.5
R5691 VSS.n14024 VSS.n14023 92.5
R5692 VSS.t32 VSS.n14037 92.5
R5693 VSS.n13907 VSS.n13906 92.5
R5694 VSS.n13894 VSS.n13893 92.5
R5695 VSS.n13859 VSS.n13858 92.5
R5696 VSS.n13853 VSS.n13852 92.5
R5697 VSS.n13855 VSS.n13854 92.5
R5698 VSS.n13848 VSS.n13847 92.5
R5699 VSS.n13850 VSS.n13849 92.5
R5700 VSS.n13844 VSS.n13843 92.5
R5701 VSS.t46 VSS.n13857 92.5
R5702 VSS.n13727 VSS.n13726 92.5
R5703 VSS.n13714 VSS.n13713 92.5
R5704 VSS.n13679 VSS.n13678 92.5
R5705 VSS.n13673 VSS.n13672 92.5
R5706 VSS.n13675 VSS.n13674 92.5
R5707 VSS.n13668 VSS.n13667 92.5
R5708 VSS.n13670 VSS.n13669 92.5
R5709 VSS.n13664 VSS.n13663 92.5
R5710 VSS.t44 VSS.n13677 92.5
R5711 VSS.n13547 VSS.n13546 92.5
R5712 VSS.n13534 VSS.n13533 92.5
R5713 VSS.n13499 VSS.n13498 92.5
R5714 VSS.n13493 VSS.n13492 92.5
R5715 VSS.n13495 VSS.n13494 92.5
R5716 VSS.n13488 VSS.n13487 92.5
R5717 VSS.n13490 VSS.n13489 92.5
R5718 VSS.n13484 VSS.n13483 92.5
R5719 VSS.t36 VSS.n13497 92.5
R5720 VSS.n13367 VSS.n13366 92.5
R5721 VSS.n13354 VSS.n13353 92.5
R5722 VSS.n13319 VSS.n13318 92.5
R5723 VSS.n13313 VSS.n13312 92.5
R5724 VSS.n13315 VSS.n13314 92.5
R5725 VSS.n13308 VSS.n13307 92.5
R5726 VSS.n13310 VSS.n13309 92.5
R5727 VSS.n13304 VSS.n13303 92.5
R5728 VSS.t34 VSS.n13317 92.5
R5729 VSS.n13187 VSS.n13186 92.5
R5730 VSS.n13174 VSS.n13173 92.5
R5731 VSS.n13139 VSS.n13138 92.5
R5732 VSS.n13133 VSS.n13132 92.5
R5733 VSS.n13135 VSS.n13134 92.5
R5734 VSS.n13128 VSS.n13127 92.5
R5735 VSS.n13130 VSS.n13129 92.5
R5736 VSS.n13124 VSS.n13123 92.5
R5737 VSS.t38 VSS.n13137 92.5
R5738 VSS.n13007 VSS.n13006 92.5
R5739 VSS.n12994 VSS.n12993 92.5
R5740 VSS.n12959 VSS.n12958 92.5
R5741 VSS.n12953 VSS.n12952 92.5
R5742 VSS.n12955 VSS.n12954 92.5
R5743 VSS.n12948 VSS.n12947 92.5
R5744 VSS.n12950 VSS.n12949 92.5
R5745 VSS.n12944 VSS.n12943 92.5
R5746 VSS.t42 VSS.n12957 92.5
R5747 VSS.n12827 VSS.n12826 92.5
R5748 VSS.n12814 VSS.n12813 92.5
R5749 VSS.n12779 VSS.n12778 92.5
R5750 VSS.n12773 VSS.n12772 92.5
R5751 VSS.n12775 VSS.n12774 92.5
R5752 VSS.n12768 VSS.n12767 92.5
R5753 VSS.n12770 VSS.n12769 92.5
R5754 VSS.n12764 VSS.n12763 92.5
R5755 VSS.t40 VSS.n12777 92.5
R5756 VSS.n12648 VSS.n12647 92.5
R5757 VSS.n9218 VSS.n9217 92.5
R5758 VSS.n9350 VSS.n9349 92.5
R5759 VSS.n9344 VSS.n9343 92.5
R5760 VSS.n9346 VSS.n9345 92.5
R5761 VSS.n9339 VSS.n9338 92.5
R5762 VSS.n9341 VSS.n9340 92.5
R5763 VSS.n9335 VSS.n9334 92.5
R5764 VSS.t48 VSS.n9348 92.5
R5765 VSS.n7167 VSS.n7166 92.5
R5766 VSS.n9386 VSS.n9385 92.5
R5767 VSS.n9518 VSS.n9517 92.5
R5768 VSS.n9512 VSS.n9511 92.5
R5769 VSS.n9514 VSS.n9513 92.5
R5770 VSS.n9507 VSS.n9506 92.5
R5771 VSS.n9509 VSS.n9508 92.5
R5772 VSS.n9503 VSS.n9502 92.5
R5773 VSS.t62 VSS.n9516 92.5
R5774 VSS.n7155 VSS.n7154 92.5
R5775 VSS.n9554 VSS.n9553 92.5
R5776 VSS.n9686 VSS.n9685 92.5
R5777 VSS.n9680 VSS.n9679 92.5
R5778 VSS.n9682 VSS.n9681 92.5
R5779 VSS.n9675 VSS.n9674 92.5
R5780 VSS.n9677 VSS.n9676 92.5
R5781 VSS.n9671 VSS.n9670 92.5
R5782 VSS.t60 VSS.n9684 92.5
R5783 VSS.n7143 VSS.n7142 92.5
R5784 VSS.n9722 VSS.n9721 92.5
R5785 VSS.n9854 VSS.n9853 92.5
R5786 VSS.n9848 VSS.n9847 92.5
R5787 VSS.n9850 VSS.n9849 92.5
R5788 VSS.n9843 VSS.n9842 92.5
R5789 VSS.n9845 VSS.n9844 92.5
R5790 VSS.n9839 VSS.n9838 92.5
R5791 VSS.t52 VSS.n9852 92.5
R5792 VSS.n7131 VSS.n7130 92.5
R5793 VSS.n9890 VSS.n9889 92.5
R5794 VSS.n10022 VSS.n10021 92.5
R5795 VSS.n10016 VSS.n10015 92.5
R5796 VSS.n10018 VSS.n10017 92.5
R5797 VSS.n10011 VSS.n10010 92.5
R5798 VSS.n10013 VSS.n10012 92.5
R5799 VSS.n10007 VSS.n10006 92.5
R5800 VSS.t50 VSS.n10020 92.5
R5801 VSS.n7119 VSS.n7118 92.5
R5802 VSS.n10058 VSS.n10057 92.5
R5803 VSS.n10190 VSS.n10189 92.5
R5804 VSS.n10184 VSS.n10183 92.5
R5805 VSS.n10186 VSS.n10185 92.5
R5806 VSS.n10179 VSS.n10178 92.5
R5807 VSS.n10181 VSS.n10180 92.5
R5808 VSS.n10175 VSS.n10174 92.5
R5809 VSS.t54 VSS.n10188 92.5
R5810 VSS.n7107 VSS.n7106 92.5
R5811 VSS.n10226 VSS.n10225 92.5
R5812 VSS.n10358 VSS.n10357 92.5
R5813 VSS.n10352 VSS.n10351 92.5
R5814 VSS.n10354 VSS.n10353 92.5
R5815 VSS.n10347 VSS.n10346 92.5
R5816 VSS.n10349 VSS.n10348 92.5
R5817 VSS.n10343 VSS.n10342 92.5
R5818 VSS.t58 VSS.n10356 92.5
R5819 VSS.n7095 VSS.n7094 92.5
R5820 VSS.n10509 VSS.n10508 92.5
R5821 VSS.n10511 VSS.n10510 92.5
R5822 VSS.n10504 VSS.n10503 92.5
R5823 VSS.n10506 VSS.n10505 92.5
R5824 VSS.n10500 VSS.n10499 92.5
R5825 VSS.t56 VSS.n10498 92.5
R5826 VSS.n2340 VSS.n2339 92.5
R5827 VSS.n2289 VSS.n2287 92.5
R5828 VSS.n2328 VSS.n2327 92.5
R5829 VSS.n2330 VSS.n2329 92.5
R5830 VSS.n2332 VSS.n2331 92.5
R5831 VSS.n2334 VSS.n2333 92.5
R5832 VSS.n2336 VSS.n2335 92.5
R5833 VSS.n2338 VSS.n2337 92.5
R5834 VSS.n2461 VSS.n2460 92.5
R5835 VSS.n2460 VSS.t24 92.5
R5836 VSS.n2355 VSS.n2354 92.5
R5837 VSS.n2353 VSS.n2352 92.5
R5838 VSS.n2351 VSS.n2350 92.5
R5839 VSS.n2349 VSS.n2348 92.5
R5840 VSS.n2347 VSS.n2346 92.5
R5841 VSS.n2345 VSS.n2344 92.5
R5842 VSS.n2343 VSS.n2342 92.5
R5843 VSS.n2341 VSS.n2298 92.5
R5844 VSS.t24 VSS.n2298 92.5
R5845 VSS.n2357 VSS.n2356 92.5
R5846 VSS.n2359 VSS.n2358 92.5
R5847 VSS.n2361 VSS.n2360 92.5
R5848 VSS.n2363 VSS.n2362 92.5
R5849 VSS.n2365 VSS.n2364 92.5
R5850 VSS.n2367 VSS.n2366 92.5
R5851 VSS.n2369 VSS.n2368 92.5
R5852 VSS.n2371 VSS.n2370 92.5
R5853 VSS.n2373 VSS.n2372 92.5
R5854 VSS.n2374 VSS.n2290 92.5
R5855 VSS.t24 VSS.n2290 92.5
R5856 VSS.n2407 VSS.n2406 92.5
R5857 VSS.n2378 VSS.n2309 92.5
R5858 VSS.n2454 VSS.n2306 92.5
R5859 VSS.n2445 VSS.n2310 92.5
R5860 VSS.n2388 VSS.n2305 92.5
R5861 VSS.n2392 VSS.n2311 92.5
R5862 VSS.n2396 VSS.n2304 92.5
R5863 VSS.n2459 VSS.n2314 92.5
R5864 VSS.n2402 VSS.n2308 92.5
R5865 VSS.n2250 VSS.n2249 92.5
R5866 VSS.n2199 VSS.n2197 92.5
R5867 VSS.n2238 VSS.n2237 92.5
R5868 VSS.n2240 VSS.n2239 92.5
R5869 VSS.n2242 VSS.n2241 92.5
R5870 VSS.n2244 VSS.n2243 92.5
R5871 VSS.n2246 VSS.n2245 92.5
R5872 VSS.n2248 VSS.n2247 92.5
R5873 VSS.n2551 VSS.n2550 92.5
R5874 VSS.n2550 VSS.t26 92.5
R5875 VSS.n2265 VSS.n2264 92.5
R5876 VSS.n2263 VSS.n2262 92.5
R5877 VSS.n2261 VSS.n2260 92.5
R5878 VSS.n2259 VSS.n2258 92.5
R5879 VSS.n2257 VSS.n2256 92.5
R5880 VSS.n2255 VSS.n2254 92.5
R5881 VSS.n2253 VSS.n2252 92.5
R5882 VSS.n2251 VSS.n2208 92.5
R5883 VSS.t26 VSS.n2208 92.5
R5884 VSS.n2267 VSS.n2266 92.5
R5885 VSS.n2269 VSS.n2268 92.5
R5886 VSS.n2271 VSS.n2270 92.5
R5887 VSS.n2273 VSS.n2272 92.5
R5888 VSS.n2275 VSS.n2274 92.5
R5889 VSS.n2277 VSS.n2276 92.5
R5890 VSS.n2279 VSS.n2278 92.5
R5891 VSS.n2281 VSS.n2280 92.5
R5892 VSS.n2283 VSS.n2282 92.5
R5893 VSS.n2284 VSS.n2200 92.5
R5894 VSS.t26 VSS.n2200 92.5
R5895 VSS.n2497 VSS.n2496 92.5
R5896 VSS.n2468 VSS.n2219 92.5
R5897 VSS.n2544 VSS.n2216 92.5
R5898 VSS.n2535 VSS.n2220 92.5
R5899 VSS.n2478 VSS.n2215 92.5
R5900 VSS.n2482 VSS.n2221 92.5
R5901 VSS.n2486 VSS.n2214 92.5
R5902 VSS.n2549 VSS.n2224 92.5
R5903 VSS.n2492 VSS.n2218 92.5
R5904 VSS.n2160 VSS.n2159 92.5
R5905 VSS.n2109 VSS.n2107 92.5
R5906 VSS.n2148 VSS.n2147 92.5
R5907 VSS.n2150 VSS.n2149 92.5
R5908 VSS.n2152 VSS.n2151 92.5
R5909 VSS.n2154 VSS.n2153 92.5
R5910 VSS.n2156 VSS.n2155 92.5
R5911 VSS.n2158 VSS.n2157 92.5
R5912 VSS.n2641 VSS.n2640 92.5
R5913 VSS.n2640 VSS.t22 92.5
R5914 VSS.n2175 VSS.n2174 92.5
R5915 VSS.n2173 VSS.n2172 92.5
R5916 VSS.n2171 VSS.n2170 92.5
R5917 VSS.n2169 VSS.n2168 92.5
R5918 VSS.n2167 VSS.n2166 92.5
R5919 VSS.n2165 VSS.n2164 92.5
R5920 VSS.n2163 VSS.n2162 92.5
R5921 VSS.n2161 VSS.n2118 92.5
R5922 VSS.t22 VSS.n2118 92.5
R5923 VSS.n2177 VSS.n2176 92.5
R5924 VSS.n2179 VSS.n2178 92.5
R5925 VSS.n2181 VSS.n2180 92.5
R5926 VSS.n2183 VSS.n2182 92.5
R5927 VSS.n2185 VSS.n2184 92.5
R5928 VSS.n2187 VSS.n2186 92.5
R5929 VSS.n2189 VSS.n2188 92.5
R5930 VSS.n2191 VSS.n2190 92.5
R5931 VSS.n2193 VSS.n2192 92.5
R5932 VSS.n2194 VSS.n2110 92.5
R5933 VSS.t22 VSS.n2110 92.5
R5934 VSS.n2587 VSS.n2586 92.5
R5935 VSS.n2558 VSS.n2129 92.5
R5936 VSS.n2634 VSS.n2126 92.5
R5937 VSS.n2625 VSS.n2130 92.5
R5938 VSS.n2568 VSS.n2125 92.5
R5939 VSS.n2572 VSS.n2131 92.5
R5940 VSS.n2576 VSS.n2124 92.5
R5941 VSS.n2639 VSS.n2134 92.5
R5942 VSS.n2582 VSS.n2128 92.5
R5943 VSS.n2070 VSS.n2069 92.5
R5944 VSS.n2019 VSS.n2017 92.5
R5945 VSS.n2058 VSS.n2057 92.5
R5946 VSS.n2060 VSS.n2059 92.5
R5947 VSS.n2062 VSS.n2061 92.5
R5948 VSS.n2064 VSS.n2063 92.5
R5949 VSS.n2066 VSS.n2065 92.5
R5950 VSS.n2068 VSS.n2067 92.5
R5951 VSS.n2731 VSS.n2730 92.5
R5952 VSS.n2730 VSS.t18 92.5
R5953 VSS.n2085 VSS.n2084 92.5
R5954 VSS.n2083 VSS.n2082 92.5
R5955 VSS.n2081 VSS.n2080 92.5
R5956 VSS.n2079 VSS.n2078 92.5
R5957 VSS.n2077 VSS.n2076 92.5
R5958 VSS.n2075 VSS.n2074 92.5
R5959 VSS.n2073 VSS.n2072 92.5
R5960 VSS.n2071 VSS.n2028 92.5
R5961 VSS.t18 VSS.n2028 92.5
R5962 VSS.n2087 VSS.n2086 92.5
R5963 VSS.n2089 VSS.n2088 92.5
R5964 VSS.n2091 VSS.n2090 92.5
R5965 VSS.n2093 VSS.n2092 92.5
R5966 VSS.n2095 VSS.n2094 92.5
R5967 VSS.n2097 VSS.n2096 92.5
R5968 VSS.n2099 VSS.n2098 92.5
R5969 VSS.n2101 VSS.n2100 92.5
R5970 VSS.n2103 VSS.n2102 92.5
R5971 VSS.n2104 VSS.n2020 92.5
R5972 VSS.t18 VSS.n2020 92.5
R5973 VSS.n2677 VSS.n2676 92.5
R5974 VSS.n2648 VSS.n2039 92.5
R5975 VSS.n2724 VSS.n2036 92.5
R5976 VSS.n2715 VSS.n2040 92.5
R5977 VSS.n2658 VSS.n2035 92.5
R5978 VSS.n2662 VSS.n2041 92.5
R5979 VSS.n2666 VSS.n2034 92.5
R5980 VSS.n2729 VSS.n2044 92.5
R5981 VSS.n2672 VSS.n2038 92.5
R5982 VSS.n1980 VSS.n1979 92.5
R5983 VSS.n1929 VSS.n1927 92.5
R5984 VSS.n1968 VSS.n1967 92.5
R5985 VSS.n1970 VSS.n1969 92.5
R5986 VSS.n1972 VSS.n1971 92.5
R5987 VSS.n1974 VSS.n1973 92.5
R5988 VSS.n1976 VSS.n1975 92.5
R5989 VSS.n1978 VSS.n1977 92.5
R5990 VSS.n2821 VSS.n2820 92.5
R5991 VSS.n2820 VSS.t20 92.5
R5992 VSS.n1995 VSS.n1994 92.5
R5993 VSS.n1993 VSS.n1992 92.5
R5994 VSS.n1991 VSS.n1990 92.5
R5995 VSS.n1989 VSS.n1988 92.5
R5996 VSS.n1987 VSS.n1986 92.5
R5997 VSS.n1985 VSS.n1984 92.5
R5998 VSS.n1983 VSS.n1982 92.5
R5999 VSS.n1981 VSS.n1938 92.5
R6000 VSS.t20 VSS.n1938 92.5
R6001 VSS.n1997 VSS.n1996 92.5
R6002 VSS.n1999 VSS.n1998 92.5
R6003 VSS.n2001 VSS.n2000 92.5
R6004 VSS.n2003 VSS.n2002 92.5
R6005 VSS.n2005 VSS.n2004 92.5
R6006 VSS.n2007 VSS.n2006 92.5
R6007 VSS.n2009 VSS.n2008 92.5
R6008 VSS.n2011 VSS.n2010 92.5
R6009 VSS.n2013 VSS.n2012 92.5
R6010 VSS.n2014 VSS.n1930 92.5
R6011 VSS.t20 VSS.n1930 92.5
R6012 VSS.n2767 VSS.n2766 92.5
R6013 VSS.n2738 VSS.n1949 92.5
R6014 VSS.n2814 VSS.n1946 92.5
R6015 VSS.n2805 VSS.n1950 92.5
R6016 VSS.n2748 VSS.n1945 92.5
R6017 VSS.n2752 VSS.n1951 92.5
R6018 VSS.n2756 VSS.n1944 92.5
R6019 VSS.n2819 VSS.n1954 92.5
R6020 VSS.n2762 VSS.n1948 92.5
R6021 VSS.n1890 VSS.n1889 92.5
R6022 VSS.n1839 VSS.n1837 92.5
R6023 VSS.n1878 VSS.n1877 92.5
R6024 VSS.n1880 VSS.n1879 92.5
R6025 VSS.n1882 VSS.n1881 92.5
R6026 VSS.n1884 VSS.n1883 92.5
R6027 VSS.n1886 VSS.n1885 92.5
R6028 VSS.n1888 VSS.n1887 92.5
R6029 VSS.n2911 VSS.n2910 92.5
R6030 VSS.n2910 VSS.t28 92.5
R6031 VSS.n1905 VSS.n1904 92.5
R6032 VSS.n1903 VSS.n1902 92.5
R6033 VSS.n1901 VSS.n1900 92.5
R6034 VSS.n1899 VSS.n1898 92.5
R6035 VSS.n1897 VSS.n1896 92.5
R6036 VSS.n1895 VSS.n1894 92.5
R6037 VSS.n1893 VSS.n1892 92.5
R6038 VSS.n1891 VSS.n1848 92.5
R6039 VSS.t28 VSS.n1848 92.5
R6040 VSS.n1907 VSS.n1906 92.5
R6041 VSS.n1909 VSS.n1908 92.5
R6042 VSS.n1911 VSS.n1910 92.5
R6043 VSS.n1913 VSS.n1912 92.5
R6044 VSS.n1915 VSS.n1914 92.5
R6045 VSS.n1917 VSS.n1916 92.5
R6046 VSS.n1919 VSS.n1918 92.5
R6047 VSS.n1921 VSS.n1920 92.5
R6048 VSS.n1923 VSS.n1922 92.5
R6049 VSS.n1924 VSS.n1840 92.5
R6050 VSS.t28 VSS.n1840 92.5
R6051 VSS.n2857 VSS.n2856 92.5
R6052 VSS.n2828 VSS.n1859 92.5
R6053 VSS.n2904 VSS.n1856 92.5
R6054 VSS.n2895 VSS.n1860 92.5
R6055 VSS.n2838 VSS.n1855 92.5
R6056 VSS.n2842 VSS.n1861 92.5
R6057 VSS.n2846 VSS.n1854 92.5
R6058 VSS.n2909 VSS.n1864 92.5
R6059 VSS.n2852 VSS.n1858 92.5
R6060 VSS.n1800 VSS.n1799 92.5
R6061 VSS.n1749 VSS.n1747 92.5
R6062 VSS.n1788 VSS.n1787 92.5
R6063 VSS.n1790 VSS.n1789 92.5
R6064 VSS.n1792 VSS.n1791 92.5
R6065 VSS.n1794 VSS.n1793 92.5
R6066 VSS.n1796 VSS.n1795 92.5
R6067 VSS.n1798 VSS.n1797 92.5
R6068 VSS.n3001 VSS.n3000 92.5
R6069 VSS.n3000 VSS.t30 92.5
R6070 VSS.n1815 VSS.n1814 92.5
R6071 VSS.n1813 VSS.n1812 92.5
R6072 VSS.n1811 VSS.n1810 92.5
R6073 VSS.n1809 VSS.n1808 92.5
R6074 VSS.n1807 VSS.n1806 92.5
R6075 VSS.n1805 VSS.n1804 92.5
R6076 VSS.n1803 VSS.n1802 92.5
R6077 VSS.n1801 VSS.n1758 92.5
R6078 VSS.t30 VSS.n1758 92.5
R6079 VSS.n1817 VSS.n1816 92.5
R6080 VSS.n1819 VSS.n1818 92.5
R6081 VSS.n1821 VSS.n1820 92.5
R6082 VSS.n1823 VSS.n1822 92.5
R6083 VSS.n1825 VSS.n1824 92.5
R6084 VSS.n1827 VSS.n1826 92.5
R6085 VSS.n1829 VSS.n1828 92.5
R6086 VSS.n1831 VSS.n1830 92.5
R6087 VSS.n1833 VSS.n1832 92.5
R6088 VSS.n1834 VSS.n1750 92.5
R6089 VSS.t30 VSS.n1750 92.5
R6090 VSS.n2947 VSS.n2946 92.5
R6091 VSS.n2918 VSS.n1769 92.5
R6092 VSS.n2994 VSS.n1766 92.5
R6093 VSS.n2985 VSS.n1770 92.5
R6094 VSS.n2928 VSS.n1765 92.5
R6095 VSS.n2932 VSS.n1771 92.5
R6096 VSS.n2936 VSS.n1764 92.5
R6097 VSS.n2999 VSS.n1774 92.5
R6098 VSS.n2942 VSS.n1768 92.5
R6099 VSS.n1710 VSS.n1709 92.5
R6100 VSS.n1659 VSS.n1657 92.5
R6101 VSS.n1698 VSS.n1697 92.5
R6102 VSS.n1700 VSS.n1699 92.5
R6103 VSS.n1702 VSS.n1701 92.5
R6104 VSS.n1704 VSS.n1703 92.5
R6105 VSS.n1706 VSS.n1705 92.5
R6106 VSS.n1708 VSS.n1707 92.5
R6107 VSS.n3091 VSS.n3090 92.5
R6108 VSS.n3090 VSS.t16 92.5
R6109 VSS.n1725 VSS.n1724 92.5
R6110 VSS.n1723 VSS.n1722 92.5
R6111 VSS.n1721 VSS.n1720 92.5
R6112 VSS.n1719 VSS.n1718 92.5
R6113 VSS.n1717 VSS.n1716 92.5
R6114 VSS.n1715 VSS.n1714 92.5
R6115 VSS.n1713 VSS.n1712 92.5
R6116 VSS.n1711 VSS.n1668 92.5
R6117 VSS.t16 VSS.n1668 92.5
R6118 VSS.n1727 VSS.n1726 92.5
R6119 VSS.n1729 VSS.n1728 92.5
R6120 VSS.n1731 VSS.n1730 92.5
R6121 VSS.n1733 VSS.n1732 92.5
R6122 VSS.n1735 VSS.n1734 92.5
R6123 VSS.n1737 VSS.n1736 92.5
R6124 VSS.n1739 VSS.n1738 92.5
R6125 VSS.n1741 VSS.n1740 92.5
R6126 VSS.n1743 VSS.n1742 92.5
R6127 VSS.n1744 VSS.n1660 92.5
R6128 VSS.t16 VSS.n1660 92.5
R6129 VSS.n3037 VSS.n3036 92.5
R6130 VSS.n3008 VSS.n1679 92.5
R6131 VSS.n3084 VSS.n1676 92.5
R6132 VSS.n3075 VSS.n1680 92.5
R6133 VSS.n3018 VSS.n1675 92.5
R6134 VSS.n3022 VSS.n1681 92.5
R6135 VSS.n3026 VSS.n1674 92.5
R6136 VSS.n3089 VSS.n1684 92.5
R6137 VSS.n3032 VSS.n1678 92.5
R6138 VSS.n6224 VSS.n6223 92.5
R6139 VSS.n6238 VSS.n6237 92.5
R6140 VSS.n6236 VSS.n6235 92.5
R6141 VSS.n6234 VSS.n6233 92.5
R6142 VSS.n6232 VSS.n6231 92.5
R6143 VSS.n6230 VSS.n6229 92.5
R6144 VSS.n6228 VSS.n6227 92.5
R6145 VSS.n6226 VSS.n6225 92.5
R6146 VSS.n6239 VSS.n6108 92.5
R6147 VSS.n6208 VSS.n6207 92.5
R6148 VSS.n6210 VSS.n6209 92.5
R6149 VSS.n6212 VSS.n6211 92.5
R6150 VSS.n6214 VSS.n6213 92.5
R6151 VSS.n6216 VSS.n6215 92.5
R6152 VSS.n6218 VSS.n6217 92.5
R6153 VSS.n6220 VSS.n6219 92.5
R6154 VSS.n6222 VSS.n6221 92.5
R6155 VSS.n6206 VSS.n6205 92.5
R6156 VSS.n6076 VSS.n6074 92.5
R6157 VSS.n6191 VSS.n6190 92.5
R6158 VSS.n6193 VSS.n6192 92.5
R6159 VSS.n6195 VSS.n6194 92.5
R6160 VSS.n6197 VSS.n6196 92.5
R6161 VSS.n6199 VSS.n6198 92.5
R6162 VSS.n6201 VSS.n6200 92.5
R6163 VSS.n6203 VSS.n6202 92.5
R6164 VSS.n6204 VSS.n6085 92.5
R6165 VSS.t64 VSS.n6085 92.5
R6166 VSS.n6077 VSS.n6075 92.5
R6167 VSS.n6124 VSS.n6081 92.5
R6168 VSS.t64 VSS.n6081 92.5
R6169 VSS.n6122 VSS.n6080 92.5
R6170 VSS.t64 VSS.n6080 92.5
R6171 VSS.n6120 VSS.n6082 92.5
R6172 VSS.t64 VSS.n6082 92.5
R6173 VSS.n6118 VSS.n6079 92.5
R6174 VSS.t64 VSS.n6079 92.5
R6175 VSS.n6116 VSS.n6083 92.5
R6176 VSS.t64 VSS.n6083 92.5
R6177 VSS.n6114 VSS.n6078 92.5
R6178 VSS.t64 VSS.n6078 92.5
R6179 VSS.n6112 VSS.n6084 92.5
R6180 VSS.t64 VSS.n6084 92.5
R6181 VSS.n6109 VSS.n6107 92.5
R6182 VSS.n6288 VSS.n6287 92.5
R6183 VSS.n6302 VSS.n6301 92.5
R6184 VSS.n6300 VSS.n6299 92.5
R6185 VSS.n6298 VSS.n6297 92.5
R6186 VSS.n6296 VSS.n6295 92.5
R6187 VSS.n6294 VSS.n6293 92.5
R6188 VSS.n6292 VSS.n6291 92.5
R6189 VSS.n6290 VSS.n6289 92.5
R6190 VSS.n6303 VSS.n5992 92.5
R6191 VSS.n6272 VSS.n6271 92.5
R6192 VSS.n6274 VSS.n6273 92.5
R6193 VSS.n6276 VSS.n6275 92.5
R6194 VSS.n6278 VSS.n6277 92.5
R6195 VSS.n6280 VSS.n6279 92.5
R6196 VSS.n6282 VSS.n6281 92.5
R6197 VSS.n6284 VSS.n6283 92.5
R6198 VSS.n6286 VSS.n6285 92.5
R6199 VSS.n6270 VSS.n6269 92.5
R6200 VSS.n5960 VSS.n5958 92.5
R6201 VSS.n6255 VSS.n6254 92.5
R6202 VSS.n6257 VSS.n6256 92.5
R6203 VSS.n6259 VSS.n6258 92.5
R6204 VSS.n6261 VSS.n6260 92.5
R6205 VSS.n6263 VSS.n6262 92.5
R6206 VSS.n6265 VSS.n6264 92.5
R6207 VSS.n6267 VSS.n6266 92.5
R6208 VSS.n6268 VSS.n5969 92.5
R6209 VSS.t76 VSS.n5969 92.5
R6210 VSS.n5961 VSS.n5959 92.5
R6211 VSS.n6008 VSS.n5965 92.5
R6212 VSS.t76 VSS.n5965 92.5
R6213 VSS.n6006 VSS.n5964 92.5
R6214 VSS.t76 VSS.n5964 92.5
R6215 VSS.n6004 VSS.n5966 92.5
R6216 VSS.t76 VSS.n5966 92.5
R6217 VSS.n6002 VSS.n5963 92.5
R6218 VSS.t76 VSS.n5963 92.5
R6219 VSS.n6000 VSS.n5967 92.5
R6220 VSS.t76 VSS.n5967 92.5
R6221 VSS.n5998 VSS.n5962 92.5
R6222 VSS.t76 VSS.n5962 92.5
R6223 VSS.n5996 VSS.n5968 92.5
R6224 VSS.t76 VSS.n5968 92.5
R6225 VSS.n5993 VSS.n5991 92.5
R6226 VSS.n6352 VSS.n6351 92.5
R6227 VSS.n6366 VSS.n6365 92.5
R6228 VSS.n6364 VSS.n6363 92.5
R6229 VSS.n6362 VSS.n6361 92.5
R6230 VSS.n6360 VSS.n6359 92.5
R6231 VSS.n6358 VSS.n6357 92.5
R6232 VSS.n6356 VSS.n6355 92.5
R6233 VSS.n6354 VSS.n6353 92.5
R6234 VSS.n6367 VSS.n5876 92.5
R6235 VSS.n6336 VSS.n6335 92.5
R6236 VSS.n6338 VSS.n6337 92.5
R6237 VSS.n6340 VSS.n6339 92.5
R6238 VSS.n6342 VSS.n6341 92.5
R6239 VSS.n6344 VSS.n6343 92.5
R6240 VSS.n6346 VSS.n6345 92.5
R6241 VSS.n6348 VSS.n6347 92.5
R6242 VSS.n6350 VSS.n6349 92.5
R6243 VSS.n6334 VSS.n6333 92.5
R6244 VSS.n5844 VSS.n5842 92.5
R6245 VSS.n6319 VSS.n6318 92.5
R6246 VSS.n6321 VSS.n6320 92.5
R6247 VSS.n6323 VSS.n6322 92.5
R6248 VSS.n6325 VSS.n6324 92.5
R6249 VSS.n6327 VSS.n6326 92.5
R6250 VSS.n6329 VSS.n6328 92.5
R6251 VSS.n6331 VSS.n6330 92.5
R6252 VSS.n6332 VSS.n5853 92.5
R6253 VSS.t74 VSS.n5853 92.5
R6254 VSS.n5845 VSS.n5843 92.5
R6255 VSS.n5892 VSS.n5849 92.5
R6256 VSS.t74 VSS.n5849 92.5
R6257 VSS.n5890 VSS.n5848 92.5
R6258 VSS.t74 VSS.n5848 92.5
R6259 VSS.n5888 VSS.n5850 92.5
R6260 VSS.t74 VSS.n5850 92.5
R6261 VSS.n5886 VSS.n5847 92.5
R6262 VSS.t74 VSS.n5847 92.5
R6263 VSS.n5884 VSS.n5851 92.5
R6264 VSS.t74 VSS.n5851 92.5
R6265 VSS.n5882 VSS.n5846 92.5
R6266 VSS.t74 VSS.n5846 92.5
R6267 VSS.n5880 VSS.n5852 92.5
R6268 VSS.t74 VSS.n5852 92.5
R6269 VSS.n5877 VSS.n5875 92.5
R6270 VSS.n6979 VSS.n6388 92.5
R6271 VSS.n6991 VSS.n6990 92.5
R6272 VSS.n6989 VSS.n6384 92.5
R6273 VSS.n6988 VSS.n6987 92.5
R6274 VSS.n6986 VSS.n6385 92.5
R6275 VSS.n6984 VSS.n6983 92.5
R6276 VSS.n6982 VSS.n6387 92.5
R6277 VSS.n6981 VSS.n6980 92.5
R6278 VSS.n6993 VSS.n6383 92.5
R6279 VSS.n6963 VSS.n6393 92.5
R6280 VSS.n6966 VSS.n6965 92.5
R6281 VSS.n6967 VSS.n6392 92.5
R6282 VSS.n6969 VSS.n6968 92.5
R6283 VSS.n6971 VSS.n6391 92.5
R6284 VSS.n6974 VSS.n6973 92.5
R6285 VSS.n6975 VSS.n6390 92.5
R6286 VSS.n6977 VSS.n6976 92.5
R6287 VSS.n6961 VSS.n6960 92.5
R6288 VSS.n6945 VSS.n6944 92.5
R6289 VSS.n6946 VSS.n6398 92.5
R6290 VSS.n6948 VSS.n6947 92.5
R6291 VSS.n6950 VSS.n6397 92.5
R6292 VSS.n6952 VSS.n6951 92.5
R6293 VSS.n6954 VSS.n6953 92.5
R6294 VSS.n6955 VSS.n6395 92.5
R6295 VSS.n6958 VSS.n6957 92.5
R6296 VSS.n6959 VSS.n6394 92.5
R6297 VSS.n6394 VSS.t68 92.5
R6298 VSS.n5789 VSS.n5787 92.5
R6299 VSS.n7038 VSS.n5790 92.5
R6300 VSS.n5790 VSS.t68 92.5
R6301 VSS.n7032 VSS.n5795 92.5
R6302 VSS.n5795 VSS.t68 92.5
R6303 VSS.n7026 VSS.n5801 92.5
R6304 VSS.n5801 VSS.t68 92.5
R6305 VSS.n7020 VSS.n5807 92.5
R6306 VSS.n5807 VSS.t68 92.5
R6307 VSS.n7014 VSS.n5813 92.5
R6308 VSS.n5813 VSS.t68 92.5
R6309 VSS.n7008 VSS.n5818 92.5
R6310 VSS.n5818 VSS.t68 92.5
R6311 VSS.n7002 VSS.n5825 92.5
R6312 VSS.n5825 VSS.t68 92.5
R6313 VSS.n6996 VSS.n5831 92.5
R6314 VSS.n6454 VSS.n6453 92.5
R6315 VSS.n6403 VSS.n6401 92.5
R6316 VSS.n6442 VSS.n6441 92.5
R6317 VSS.n6444 VSS.n6443 92.5
R6318 VSS.n6446 VSS.n6445 92.5
R6319 VSS.n6448 VSS.n6447 92.5
R6320 VSS.n6450 VSS.n6449 92.5
R6321 VSS.n6452 VSS.n6451 92.5
R6322 VSS.n6935 VSS.n6934 92.5
R6323 VSS.n6934 VSS.t66 92.5
R6324 VSS.n6469 VSS.n6468 92.5
R6325 VSS.n6467 VSS.n6466 92.5
R6326 VSS.n6465 VSS.n6464 92.5
R6327 VSS.n6463 VSS.n6462 92.5
R6328 VSS.n6461 VSS.n6460 92.5
R6329 VSS.n6459 VSS.n6458 92.5
R6330 VSS.n6457 VSS.n6456 92.5
R6331 VSS.n6455 VSS.n6412 92.5
R6332 VSS.t66 VSS.n6412 92.5
R6333 VSS.n6471 VSS.n6470 92.5
R6334 VSS.n6473 VSS.n6472 92.5
R6335 VSS.n6475 VSS.n6474 92.5
R6336 VSS.n6477 VSS.n6476 92.5
R6337 VSS.n6479 VSS.n6478 92.5
R6338 VSS.n6481 VSS.n6480 92.5
R6339 VSS.n6483 VSS.n6482 92.5
R6340 VSS.n6485 VSS.n6484 92.5
R6341 VSS.n6487 VSS.n6486 92.5
R6342 VSS.n6488 VSS.n6404 92.5
R6343 VSS.t66 VSS.n6404 92.5
R6344 VSS.n6852 VSS.n6851 92.5
R6345 VSS.n6927 VSS.n6423 92.5
R6346 VSS.n6918 VSS.n6420 92.5
R6347 VSS.n6862 VSS.n6424 92.5
R6348 VSS.n6866 VSS.n6419 92.5
R6349 VSS.n6870 VSS.n6425 92.5
R6350 VSS.n6874 VSS.n6418 92.5
R6351 VSS.n6933 VSS.n6428 92.5
R6352 VSS.n6880 VSS.n6422 92.5
R6353 VSS.n6544 VSS.n6543 92.5
R6354 VSS.n6493 VSS.n6491 92.5
R6355 VSS.n6532 VSS.n6531 92.5
R6356 VSS.n6534 VSS.n6533 92.5
R6357 VSS.n6536 VSS.n6535 92.5
R6358 VSS.n6538 VSS.n6537 92.5
R6359 VSS.n6540 VSS.n6539 92.5
R6360 VSS.n6542 VSS.n6541 92.5
R6361 VSS.n6845 VSS.n6844 92.5
R6362 VSS.n6844 VSS.t70 92.5
R6363 VSS.n6559 VSS.n6558 92.5
R6364 VSS.n6557 VSS.n6556 92.5
R6365 VSS.n6555 VSS.n6554 92.5
R6366 VSS.n6553 VSS.n6552 92.5
R6367 VSS.n6551 VSS.n6550 92.5
R6368 VSS.n6549 VSS.n6548 92.5
R6369 VSS.n6547 VSS.n6546 92.5
R6370 VSS.n6545 VSS.n6502 92.5
R6371 VSS.t70 VSS.n6502 92.5
R6372 VSS.n6561 VSS.n6560 92.5
R6373 VSS.n6563 VSS.n6562 92.5
R6374 VSS.n6565 VSS.n6564 92.5
R6375 VSS.n6567 VSS.n6566 92.5
R6376 VSS.n6569 VSS.n6568 92.5
R6377 VSS.n6571 VSS.n6570 92.5
R6378 VSS.n6573 VSS.n6572 92.5
R6379 VSS.n6575 VSS.n6574 92.5
R6380 VSS.n6577 VSS.n6576 92.5
R6381 VSS.n6578 VSS.n6494 92.5
R6382 VSS.t70 VSS.n6494 92.5
R6383 VSS.n6762 VSS.n6761 92.5
R6384 VSS.n6837 VSS.n6513 92.5
R6385 VSS.n6828 VSS.n6510 92.5
R6386 VSS.n6772 VSS.n6514 92.5
R6387 VSS.n6776 VSS.n6509 92.5
R6388 VSS.n6780 VSS.n6515 92.5
R6389 VSS.n6784 VSS.n6508 92.5
R6390 VSS.n6843 VSS.n6518 92.5
R6391 VSS.n6790 VSS.n6512 92.5
R6392 VSS.n6634 VSS.n6633 92.5
R6393 VSS.n6583 VSS.n6581 92.5
R6394 VSS.n6622 VSS.n6621 92.5
R6395 VSS.n6624 VSS.n6623 92.5
R6396 VSS.n6626 VSS.n6625 92.5
R6397 VSS.n6628 VSS.n6627 92.5
R6398 VSS.n6630 VSS.n6629 92.5
R6399 VSS.n6632 VSS.n6631 92.5
R6400 VSS.n6755 VSS.n6754 92.5
R6401 VSS.n6754 VSS.t72 92.5
R6402 VSS.n6649 VSS.n6648 92.5
R6403 VSS.n6647 VSS.n6646 92.5
R6404 VSS.n6645 VSS.n6644 92.5
R6405 VSS.n6643 VSS.n6642 92.5
R6406 VSS.n6641 VSS.n6640 92.5
R6407 VSS.n6639 VSS.n6638 92.5
R6408 VSS.n6637 VSS.n6636 92.5
R6409 VSS.n6635 VSS.n6592 92.5
R6410 VSS.t72 VSS.n6592 92.5
R6411 VSS.n6651 VSS.n6650 92.5
R6412 VSS.n6653 VSS.n6652 92.5
R6413 VSS.n6655 VSS.n6654 92.5
R6414 VSS.n6657 VSS.n6656 92.5
R6415 VSS.n6659 VSS.n6658 92.5
R6416 VSS.n6661 VSS.n6660 92.5
R6417 VSS.n6663 VSS.n6662 92.5
R6418 VSS.n6665 VSS.n6664 92.5
R6419 VSS.n6667 VSS.n6666 92.5
R6420 VSS.n6668 VSS.n6584 92.5
R6421 VSS.t72 VSS.n6584 92.5
R6422 VSS.n6672 VSS.n6671 92.5
R6423 VSS.n6747 VSS.n6603 92.5
R6424 VSS.n6738 VSS.n6600 92.5
R6425 VSS.n6682 VSS.n6604 92.5
R6426 VSS.n6686 VSS.n6599 92.5
R6427 VSS.n6690 VSS.n6605 92.5
R6428 VSS.n6694 VSS.n6598 92.5
R6429 VSS.n6753 VSS.n6608 92.5
R6430 VSS.n6700 VSS.n6602 92.5
R6431 VSS.n17998 VSS.n17997 92.5
R6432 VSS.n18012 VSS.n18011 92.5
R6433 VSS.n18010 VSS.n18009 92.5
R6434 VSS.n18008 VSS.n18007 92.5
R6435 VSS.n18006 VSS.n18005 92.5
R6436 VSS.n18004 VSS.n18003 92.5
R6437 VSS.n18002 VSS.n18001 92.5
R6438 VSS.n18000 VSS.n17999 92.5
R6439 VSS.n18013 VSS.n17946 92.5
R6440 VSS.n17996 VSS.n17995 92.5
R6441 VSS.n17994 VSS.n17993 92.5
R6442 VSS.n17992 VSS.n17991 92.5
R6443 VSS.n17990 VSS.n17989 92.5
R6444 VSS.n17988 VSS.n17987 92.5
R6445 VSS.n17986 VSS.n17985 92.5
R6446 VSS.n17984 VSS.n17983 92.5
R6447 VSS.n17982 VSS.n17981 92.5
R6448 VSS.n17980 VSS.n17979 92.5
R6449 VSS.n17978 VSS.n17977 92.5
R6450 VSS.n17976 VSS.n17975 92.5
R6451 VSS.n17974 VSS.n17973 92.5
R6452 VSS.n17972 VSS.n17971 92.5
R6453 VSS.n17970 VSS.n17969 92.5
R6454 VSS.n17968 VSS.n17967 92.5
R6455 VSS.n17966 VSS.n17965 92.5
R6456 VSS.n17964 VSS.n17963 92.5
R6457 VSS.n17962 VSS.n17961 92.5
R6458 VSS.n17950 VSS.n17949 92.5
R6459 VSS.n17952 VSS.n17951 92.5
R6460 VSS.n17954 VSS.n17953 92.5
R6461 VSS.n17956 VSS.n17955 92.5
R6462 VSS.n17958 VSS.n17957 92.5
R6463 VSS.n17960 VSS.n17959 92.5
R6464 VSS.n18015 VSS.n18014 92.5
R6465 VSS.n17947 VSS.n17922 92.5
R6466 VSS.n497 VSS.n471 91.028
R6467 VSS.n15107 VSS.n15106 89.722
R6468 VSS.n14862 VSS.n14861 89.722
R6469 VSS.n15595 VSS.n15594 89.722
R6470 VSS.n15350 VSS.n15349 89.722
R6471 VSS.n16083 VSS.n16082 89.722
R6472 VSS.n15838 VSS.n15837 89.722
R6473 VSS.n16338 VSS.n16337 89.722
R6474 VSS.n11156 VSS.n11155 89.722
R6475 VSS.n10911 VSS.n10910 89.722
R6476 VSS.n11644 VSS.n11643 89.722
R6477 VSS.n11399 VSS.n11398 89.722
R6478 VSS.n12132 VSS.n12131 89.722
R6479 VSS.n11887 VSS.n11886 89.722
R6480 VSS.n12387 VSS.n12386 89.722
R6481 VSS.n7724 VSS.n7723 89.722
R6482 VSS.n7479 VSS.n7478 89.722
R6483 VSS.n8212 VSS.n8211 89.722
R6484 VSS.n7967 VSS.n7966 89.722
R6485 VSS.n8700 VSS.n8699 89.722
R6486 VSS.n8455 VSS.n8454 89.722
R6487 VSS.n8955 VSS.n8954 89.722
R6488 VSS.n5463 VSS.n1461 89.722
R6489 VSS.n5438 VSS.n1507 89.722
R6490 VSS.n5671 VSS.n606 89.722
R6491 VSS.n5646 VSS.n1366 89.722
R6492 VSS.n1299 VSS.n636 89.722
R6493 VSS.n622 VSS.n618 89.722
R6494 VSS.n3923 VSS.n3408 89.722
R6495 VSS.n3859 VSS.n3422 89.722
R6496 VSS.n4472 VSS.n3293 89.722
R6497 VSS.n3898 VSS.n3306 89.722
R6498 VSS.n3254 VSS.n3139 89.722
R6499 VSS.n4501 VSS.n3242 89.722
R6500 VSS.n5074 VSS.n3126 89.722
R6501 VSS.n2458 VSS.n2315 89.673
R6502 VSS.n2548 VSS.n2225 89.673
R6503 VSS.n2638 VSS.n2135 89.673
R6504 VSS.n2728 VSS.n2045 89.673
R6505 VSS.n2818 VSS.n1955 89.673
R6506 VSS.n2908 VSS.n1865 89.673
R6507 VSS.n2998 VSS.n1775 89.673
R6508 VSS.n3088 VSS.n1685 89.673
R6509 VSS.n5495 VSS.n1445 83.871
R6510 VSS.n5399 VSS.n1527 83.871
R6511 VSS.n781 VSS.n592 83.871
R6512 VSS.n5607 VSS.n1386 83.871
R6513 VSS.n717 VSS.n714 83.871
R6514 VSS.n1022 VSS.n651 83.871
R6515 VSS.n3388 VSS.n3384 83.871
R6516 VSS.n3565 VSS.n3523 83.871
R6517 VSS.n4177 VSS.n4135 83.871
R6518 VSS.n4064 VSS.n3321 83.871
R6519 VSS.n4655 VSS.n3154 83.871
R6520 VSS.n4530 VSS.n3217 83.871
R6521 VSS.n4767 VSS.n4725 83.871
R6522 VSS.n2457 VSS.n2456 71.237
R6523 VSS.n2446 VSS.n2316 71.237
R6524 VSS.n2386 VSS.n2322 71.237
R6525 VSS.n2389 VSS.n2317 71.237
R6526 VSS.n2393 VSS.n2321 71.237
R6527 VSS.n2320 VSS.n2312 71.237
R6528 VSS.n2399 VSS.n2319 71.237
R6529 VSS.n2405 VSS.n2318 71.237
R6530 VSS.n2547 VSS.n2546 71.237
R6531 VSS.n2536 VSS.n2226 71.237
R6532 VSS.n2476 VSS.n2232 71.237
R6533 VSS.n2479 VSS.n2227 71.237
R6534 VSS.n2483 VSS.n2231 71.237
R6535 VSS.n2230 VSS.n2222 71.237
R6536 VSS.n2489 VSS.n2229 71.237
R6537 VSS.n2495 VSS.n2228 71.237
R6538 VSS.n2637 VSS.n2636 71.237
R6539 VSS.n2626 VSS.n2136 71.237
R6540 VSS.n2566 VSS.n2142 71.237
R6541 VSS.n2569 VSS.n2137 71.237
R6542 VSS.n2573 VSS.n2141 71.237
R6543 VSS.n2140 VSS.n2132 71.237
R6544 VSS.n2579 VSS.n2139 71.237
R6545 VSS.n2585 VSS.n2138 71.237
R6546 VSS.n2727 VSS.n2726 71.237
R6547 VSS.n2716 VSS.n2046 71.237
R6548 VSS.n2656 VSS.n2052 71.237
R6549 VSS.n2659 VSS.n2047 71.237
R6550 VSS.n2663 VSS.n2051 71.237
R6551 VSS.n2050 VSS.n2042 71.237
R6552 VSS.n2669 VSS.n2049 71.237
R6553 VSS.n2675 VSS.n2048 71.237
R6554 VSS.n2817 VSS.n2816 71.237
R6555 VSS.n2806 VSS.n1956 71.237
R6556 VSS.n2746 VSS.n1962 71.237
R6557 VSS.n2749 VSS.n1957 71.237
R6558 VSS.n2753 VSS.n1961 71.237
R6559 VSS.n1960 VSS.n1952 71.237
R6560 VSS.n2759 VSS.n1959 71.237
R6561 VSS.n2765 VSS.n1958 71.237
R6562 VSS.n2907 VSS.n2906 71.237
R6563 VSS.n2896 VSS.n1866 71.237
R6564 VSS.n2836 VSS.n1872 71.237
R6565 VSS.n2839 VSS.n1867 71.237
R6566 VSS.n2843 VSS.n1871 71.237
R6567 VSS.n1870 VSS.n1862 71.237
R6568 VSS.n2849 VSS.n1869 71.237
R6569 VSS.n2855 VSS.n1868 71.237
R6570 VSS.n2997 VSS.n2996 71.237
R6571 VSS.n2986 VSS.n1776 71.237
R6572 VSS.n2926 VSS.n1782 71.237
R6573 VSS.n2929 VSS.n1777 71.237
R6574 VSS.n2933 VSS.n1781 71.237
R6575 VSS.n1780 VSS.n1772 71.237
R6576 VSS.n2939 VSS.n1779 71.237
R6577 VSS.n2945 VSS.n1778 71.237
R6578 VSS.n3087 VSS.n3086 71.237
R6579 VSS.n3076 VSS.n1686 71.237
R6580 VSS.n3016 VSS.n1692 71.237
R6581 VSS.n3019 VSS.n1687 71.237
R6582 VSS.n3023 VSS.n1691 71.237
R6583 VSS.n1690 VSS.n1682 71.237
R6584 VSS.n3029 VSS.n1689 71.237
R6585 VSS.n3035 VSS.n1688 71.237
R6586 VSS.n6129 VSS.n6105 71.237
R6587 VSS.n6137 VSS.n6104 71.237
R6588 VSS.n6145 VSS.n6100 71.237
R6589 VSS.n6153 VSS.n6101 71.237
R6590 VSS.n6161 VSS.n6106 71.237
R6591 VSS.n6169 VSS.n6103 71.237
R6592 VSS.n6177 VSS.n6099 71.237
R6593 VSS.n6185 VSS.n6102 71.237
R6594 VSS.n6013 VSS.n5989 71.237
R6595 VSS.n6021 VSS.n5988 71.237
R6596 VSS.n6029 VSS.n5984 71.237
R6597 VSS.n6037 VSS.n5985 71.237
R6598 VSS.n6045 VSS.n5990 71.237
R6599 VSS.n6053 VSS.n5987 71.237
R6600 VSS.n6061 VSS.n5983 71.237
R6601 VSS.n6069 VSS.n5986 71.237
R6602 VSS.n5897 VSS.n5873 71.237
R6603 VSS.n5905 VSS.n5872 71.237
R6604 VSS.n5913 VSS.n5868 71.237
R6605 VSS.n5921 VSS.n5869 71.237
R6606 VSS.n5929 VSS.n5874 71.237
R6607 VSS.n5937 VSS.n5871 71.237
R6608 VSS.n5945 VSS.n5867 71.237
R6609 VSS.n5953 VSS.n5870 71.237
R6610 VSS.n7041 VSS.n7040 71.237
R6611 VSS.n7035 VSS.n7034 71.237
R6612 VSS.n7029 VSS.n7028 71.237
R6613 VSS.n7023 VSS.n7022 71.237
R6614 VSS.n7017 VSS.n7016 71.237
R6615 VSS.n7011 VSS.n7010 71.237
R6616 VSS.n7005 VSS.n7004 71.237
R6617 VSS.n6999 VSS.n6998 71.237
R6618 VSS.n6930 VSS.n6929 71.237
R6619 VSS.n6919 VSS.n6430 71.237
R6620 VSS.n6860 VSS.n6436 71.237
R6621 VSS.n6863 VSS.n6431 71.237
R6622 VSS.n6867 VSS.n6435 71.237
R6623 VSS.n6871 VSS.n6432 71.237
R6624 VSS.n6434 VSS.n6426 71.237
R6625 VSS.n6877 VSS.n6433 71.237
R6626 VSS.n6840 VSS.n6839 71.237
R6627 VSS.n6829 VSS.n6520 71.237
R6628 VSS.n6770 VSS.n6526 71.237
R6629 VSS.n6773 VSS.n6521 71.237
R6630 VSS.n6777 VSS.n6525 71.237
R6631 VSS.n6781 VSS.n6522 71.237
R6632 VSS.n6524 VSS.n6516 71.237
R6633 VSS.n6787 VSS.n6523 71.237
R6634 VSS.n6750 VSS.n6749 71.237
R6635 VSS.n6739 VSS.n6610 71.237
R6636 VSS.n6680 VSS.n6616 71.237
R6637 VSS.n6683 VSS.n6611 71.237
R6638 VSS.n6687 VSS.n6615 71.237
R6639 VSS.n6691 VSS.n6612 71.237
R6640 VSS.n6614 VSS.n6606 71.237
R6641 VSS.n6697 VSS.n6613 71.237
R6642 VSS.n14807 VSS.n14802 70.217
R6643 VSS.n15307 VSS.n15302 70.217
R6644 VSS.n15063 VSS.n15058 70.217
R6645 VSS.n15795 VSS.n15790 70.217
R6646 VSS.n15551 VSS.n15546 70.217
R6647 VSS.n16283 VSS.n16278 70.217
R6648 VSS.n16039 VSS.n16034 70.217
R6649 VSS.n10856 VSS.n10851 70.217
R6650 VSS.n11356 VSS.n11351 70.217
R6651 VSS.n11112 VSS.n11107 70.217
R6652 VSS.n11844 VSS.n11839 70.217
R6653 VSS.n11600 VSS.n11595 70.217
R6654 VSS.n12332 VSS.n12327 70.217
R6655 VSS.n12088 VSS.n12083 70.217
R6656 VSS.n7424 VSS.n7419 70.217
R6657 VSS.n7924 VSS.n7919 70.217
R6658 VSS.n7680 VSS.n7675 70.217
R6659 VSS.n8412 VSS.n8407 70.217
R6660 VSS.n8168 VSS.n8163 70.217
R6661 VSS.n8900 VSS.n8895 70.217
R6662 VSS.n8656 VSS.n8651 70.217
R6663 VSS.n5403 VSS.n1527 70.217
R6664 VSS.n5611 VSS.n1386 70.217
R6665 VSS.n5310 VSS.n1445 70.217
R6666 VSS.n879 VSS.n717 70.217
R6667 VSS.n592 VSS.n584 70.217
R6668 VSS.n1267 VSS.n651 70.217
R6669 VSS.n3720 VSS.n3523 70.217
R6670 VSS.n4418 VSS.n3321 70.217
R6671 VSS.n3957 VSS.n3388 70.217
R6672 VSS.n4531 VSS.n4530 70.217
R6673 VSS.n4324 VSS.n4135 70.217
R6674 VSS.n4933 VSS.n4725 70.217
R6675 VSS.n4645 VSS.n3154 70.217
R6676 VSS.n5412 VSS.n1520 69.803
R6677 VSS.n5412 VSS.n1518 69.803
R6678 VSS.n5416 VSS.n1518 69.803
R6679 VSS.n5416 VSS.n1516 69.803
R6680 VSS.n5420 VSS.n1516 69.803
R6681 VSS.n5420 VSS.n1514 69.803
R6682 VSS.n5424 VSS.n1514 69.803
R6683 VSS.n5424 VSS.n1512 69.803
R6684 VSS.n5429 VSS.n1512 69.803
R6685 VSS.n5429 VSS.n1510 69.803
R6686 VSS.n5433 VSS.n1510 69.803
R6687 VSS.n5434 VSS.n5433 69.803
R6688 VSS.n5491 VSS.n1449 69.803
R6689 VSS.n5487 VSS.n1449 69.803
R6690 VSS.n5487 VSS.n1451 69.803
R6691 VSS.n5483 VSS.n1451 69.803
R6692 VSS.n5483 VSS.n1453 69.803
R6693 VSS.n5479 VSS.n1453 69.803
R6694 VSS.n5479 VSS.n1455 69.803
R6695 VSS.n5475 VSS.n1455 69.803
R6696 VSS.n5475 VSS.n1457 69.803
R6697 VSS.n5471 VSS.n1457 69.803
R6698 VSS.n5471 VSS.n1459 69.803
R6699 VSS.n5467 VSS.n1459 69.803
R6700 VSS.n5620 VSS.n1379 69.803
R6701 VSS.n5620 VSS.n1377 69.803
R6702 VSS.n5624 VSS.n1377 69.803
R6703 VSS.n5624 VSS.n1375 69.803
R6704 VSS.n5628 VSS.n1375 69.803
R6705 VSS.n5628 VSS.n1373 69.803
R6706 VSS.n5632 VSS.n1373 69.803
R6707 VSS.n5632 VSS.n1371 69.803
R6708 VSS.n5637 VSS.n1371 69.803
R6709 VSS.n5637 VSS.n1369 69.803
R6710 VSS.n5641 VSS.n1369 69.803
R6711 VSS.n5642 VSS.n5641 69.803
R6712 VSS.n5699 VSS.n593 69.803
R6713 VSS.n5695 VSS.n593 69.803
R6714 VSS.n5695 VSS.n596 69.803
R6715 VSS.n5691 VSS.n596 69.803
R6716 VSS.n5691 VSS.n598 69.803
R6717 VSS.n5687 VSS.n598 69.803
R6718 VSS.n5687 VSS.n600 69.803
R6719 VSS.n5683 VSS.n600 69.803
R6720 VSS.n5683 VSS.n602 69.803
R6721 VSS.n5679 VSS.n602 69.803
R6722 VSS.n5679 VSS.n604 69.803
R6723 VSS.n5675 VSS.n604 69.803
R6724 VSS.n915 VSS.n718 69.803
R6725 VSS.n911 VSS.n718 69.803
R6726 VSS.n911 VSS.n887 69.803
R6727 VSS.n907 VSS.n887 69.803
R6728 VSS.n907 VSS.n889 69.803
R6729 VSS.n903 VSS.n889 69.803
R6730 VSS.n903 VSS.n891 69.803
R6731 VSS.n899 VSS.n891 69.803
R6732 VSS.n899 VSS.n893 69.803
R6733 VSS.n895 VSS.n893 69.803
R6734 VSS.n895 VSS.n621 69.803
R6735 VSS.n1324 VSS.n621 69.803
R6736 VSS.n1271 VSS.n649 69.803
R6737 VSS.n1275 VSS.n649 69.803
R6738 VSS.n1275 VSS.n647 69.803
R6739 VSS.n1279 VSS.n647 69.803
R6740 VSS.n1279 VSS.n645 69.803
R6741 VSS.n1283 VSS.n645 69.803
R6742 VSS.n1283 VSS.n643 69.803
R6743 VSS.n1287 VSS.n643 69.803
R6744 VSS.n1287 VSS.n641 69.803
R6745 VSS.n1291 VSS.n641 69.803
R6746 VSS.n1291 VSS.n639 69.803
R6747 VSS.n1295 VSS.n639 69.803
R6748 VSS.n3556 VSS.n3526 69.803
R6749 VSS.n3552 VSS.n3526 69.803
R6750 VSS.n3552 VSS.n3528 69.803
R6751 VSS.n3548 VSS.n3528 69.803
R6752 VSS.n3548 VSS.n3530 69.803
R6753 VSS.n3544 VSS.n3530 69.803
R6754 VSS.n3544 VSS.n3532 69.803
R6755 VSS.n3540 VSS.n3532 69.803
R6756 VSS.n3540 VSS.n3534 69.803
R6757 VSS.n3536 VSS.n3534 69.803
R6758 VSS.n3536 VSS.n3421 69.803
R6759 VSS.n3863 VSS.n3421 69.803
R6760 VSS.n3949 VSS.n3948 69.803
R6761 VSS.n3948 VSS.n3393 69.803
R6762 VSS.n3944 VSS.n3393 69.803
R6763 VSS.n3944 VSS.n3395 69.803
R6764 VSS.n3940 VSS.n3395 69.803
R6765 VSS.n3940 VSS.n3398 69.803
R6766 VSS.n3936 VSS.n3398 69.803
R6767 VSS.n3936 VSS.n3400 69.803
R6768 VSS.n3932 VSS.n3400 69.803
R6769 VSS.n3932 VSS.n3402 69.803
R6770 VSS.n3928 VSS.n3402 69.803
R6771 VSS.n3928 VSS.n3404 69.803
R6772 VSS.n4422 VSS.n3319 69.803
R6773 VSS.n4426 VSS.n3319 69.803
R6774 VSS.n4426 VSS.n3317 69.803
R6775 VSS.n4430 VSS.n3317 69.803
R6776 VSS.n4430 VSS.n3315 69.803
R6777 VSS.n4434 VSS.n3315 69.803
R6778 VSS.n4434 VSS.n3313 69.803
R6779 VSS.n4438 VSS.n3313 69.803
R6780 VSS.n4438 VSS.n3311 69.803
R6781 VSS.n4442 VSS.n3311 69.803
R6782 VSS.n4442 VSS.n3309 69.803
R6783 VSS.n4446 VSS.n3309 69.803
R6784 VSS.n4168 VSS.n4138 69.803
R6785 VSS.n4164 VSS.n4138 69.803
R6786 VSS.n4164 VSS.n4140 69.803
R6787 VSS.n4160 VSS.n4140 69.803
R6788 VSS.n4160 VSS.n4142 69.803
R6789 VSS.n4156 VSS.n4142 69.803
R6790 VSS.n4156 VSS.n4144 69.803
R6791 VSS.n4152 VSS.n4144 69.803
R6792 VSS.n4152 VSS.n4146 69.803
R6793 VSS.n4148 VSS.n4146 69.803
R6794 VSS.n4148 VSS.n3292 69.803
R6795 VSS.n4476 VSS.n3292 69.803
R6796 VSS.n4529 VSS.n3229 69.803
R6797 VSS.n4525 VSS.n3229 69.803
R6798 VSS.n4525 VSS.n3231 69.803
R6799 VSS.n4521 VSS.n3231 69.803
R6800 VSS.n4521 VSS.n3234 69.803
R6801 VSS.n4517 VSS.n3234 69.803
R6802 VSS.n4517 VSS.n3236 69.803
R6803 VSS.n4513 VSS.n3236 69.803
R6804 VSS.n4513 VSS.n3238 69.803
R6805 VSS.n4509 VSS.n3238 69.803
R6806 VSS.n4509 VSS.n3240 69.803
R6807 VSS.n4505 VSS.n3240 69.803
R6808 VSS.n5024 VSS.n3152 69.803
R6809 VSS.n5028 VSS.n3152 69.803
R6810 VSS.n5028 VSS.n3150 69.803
R6811 VSS.n5032 VSS.n3150 69.803
R6812 VSS.n5032 VSS.n3148 69.803
R6813 VSS.n5036 VSS.n3148 69.803
R6814 VSS.n5036 VSS.n3146 69.803
R6815 VSS.n5040 VSS.n3146 69.803
R6816 VSS.n5040 VSS.n3144 69.803
R6817 VSS.n5044 VSS.n3144 69.803
R6818 VSS.n5044 VSS.n3142 69.803
R6819 VSS.n5048 VSS.n3142 69.803
R6820 VSS.n4758 VSS.n4728 69.803
R6821 VSS.n4754 VSS.n4728 69.803
R6822 VSS.n4754 VSS.n4730 69.803
R6823 VSS.n4750 VSS.n4730 69.803
R6824 VSS.n4750 VSS.n4732 69.803
R6825 VSS.n4746 VSS.n4732 69.803
R6826 VSS.n4746 VSS.n4734 69.803
R6827 VSS.n4742 VSS.n4734 69.803
R6828 VSS.n4742 VSS.n4736 69.803
R6829 VSS.n4738 VSS.n4736 69.803
R6830 VSS.n4738 VSS.n3125 69.803
R6831 VSS.n5078 VSS.n3125 69.803
R6832 VSS.n17997 VSS.n17938 68.545
R6833 VSS.t78 VSS.n17944 65.818
R6834 VSS.t78 VSS.n17943 65.818
R6835 VSS.t78 VSS.n17942 65.818
R6836 VSS.t78 VSS.n17941 65.818
R6837 VSS.t78 VSS.n17940 65.818
R6838 VSS.t78 VSS.n17939 65.818
R6839 VSS.n18009 VSS.n17945 64.913
R6840 VSS.n14864 VSS.n14862 64.374
R6841 VSS.n15109 VSS.n15107 64.374
R6842 VSS.n15352 VSS.n15350 64.374
R6843 VSS.n15597 VSS.n15595 64.374
R6844 VSS.n15840 VSS.n15838 64.374
R6845 VSS.n16085 VSS.n16083 64.374
R6846 VSS.n16340 VSS.n16338 64.374
R6847 VSS.n10913 VSS.n10911 64.374
R6848 VSS.n11158 VSS.n11156 64.374
R6849 VSS.n11401 VSS.n11399 64.374
R6850 VSS.n11646 VSS.n11644 64.374
R6851 VSS.n11889 VSS.n11887 64.374
R6852 VSS.n12134 VSS.n12132 64.374
R6853 VSS.n12389 VSS.n12387 64.374
R6854 VSS.n7481 VSS.n7479 64.374
R6855 VSS.n7726 VSS.n7724 64.374
R6856 VSS.n7969 VSS.n7967 64.374
R6857 VSS.n8214 VSS.n8212 64.374
R6858 VSS.n8457 VSS.n8455 64.374
R6859 VSS.n8702 VSS.n8700 64.374
R6860 VSS.n8957 VSS.n8955 64.374
R6861 VSS.n5434 VSS.n1507 64.374
R6862 VSS.n5467 VSS.n1461 64.374
R6863 VSS.n5642 VSS.n1366 64.374
R6864 VSS.n5675 VSS.n606 64.374
R6865 VSS.n1324 VSS.n622 64.374
R6866 VSS.n1295 VSS.n636 64.374
R6867 VSS.n3863 VSS.n3422 64.374
R6868 VSS.n3408 VSS.n3404 64.374
R6869 VSS.n4446 VSS.n3306 64.374
R6870 VSS.n4476 VSS.n3293 64.374
R6871 VSS.n4505 VSS.n3242 64.374
R6872 VSS.n5048 VSS.n3139 64.374
R6873 VSS.n5078 VSS.n3126 64.374
R6874 VSS.n6248 VSS.t64 59.179
R6875 VSS.n6312 VSS.t76 59.179
R6876 VSS.n6376 VSS.t74 59.179
R6877 VSS.n6941 VSS.t68 59.179
R6878 VSS.n17927 VSS.n17925 57.98
R6879 VSS.n17947 VSS.n17924 54.346
R6880 VSS.n17550 VSS.n17548 53.901
R6881 VSS.n17550 VSS.n17549 53.901
R6882 VSS.n17382 VSS.n17380 53.901
R6883 VSS.n17382 VSS.n17381 53.901
R6884 VSS.n17214 VSS.n17212 53.901
R6885 VSS.n17214 VSS.n17213 53.901
R6886 VSS.n17046 VSS.n17044 53.901
R6887 VSS.n17046 VSS.n17045 53.901
R6888 VSS.n16878 VSS.n16876 53.901
R6889 VSS.n16878 VSS.n16877 53.901
R6890 VSS.n16710 VSS.n16708 53.901
R6891 VSS.n16710 VSS.n16709 53.901
R6892 VSS.n10515 VSS.n10513 53.901
R6893 VSS.n10515 VSS.n10514 53.901
R6894 VSS.n6221 VSS.n6089 53.901
R6895 VSS.n6224 VSS.n6089 53.901
R6896 VSS.n6285 VSS.n5973 53.901
R6897 VSS.n6288 VSS.n5973 53.901
R6898 VSS.n6349 VSS.n5857 53.901
R6899 VSS.n6352 VSS.n5857 53.901
R6900 VSS.n6978 VSS.n6977 53.901
R6901 VSS.n6979 VSS.n6978 53.901
R6902 VSS.n17959 VSS.n17936 53.901
R6903 VSS.n17962 VSS.n17936 53.901
R6904 VSS.n17999 VSS.n17939 53.366
R6905 VSS.n18001 VSS.n17940 53.366
R6906 VSS.n18003 VSS.n17941 53.366
R6907 VSS.n18005 VSS.n17942 53.366
R6908 VSS.n18007 VSS.n17943 53.366
R6909 VSS.n18009 VSS.n17944 53.366
R6910 VSS.n17999 VSS.n17940 53.366
R6911 VSS.n18001 VSS.n17941 53.366
R6912 VSS.n18003 VSS.n17942 53.366
R6913 VSS.n18005 VSS.n17943 53.366
R6914 VSS.n18007 VSS.n17944 53.366
R6915 VSS.n17997 VSS.n17939 53.366
R6916 VSS.n18016 VSS.n18015 53.161
R6917 VSS.n18016 VSS.n17946 53.161
R6918 VSS.t78 VSS.n17927 42.341
R6919 VSS.n14444 VSS.n14442 41.419
R6920 VSS.n14439 VSS.n14436 41.419
R6921 VSS.n14434 VSS.n14431 41.419
R6922 VSS.n14429 VSS.n14427 41.419
R6923 VSS.n14264 VSS.n14262 41.419
R6924 VSS.n14259 VSS.n14256 41.419
R6925 VSS.n14254 VSS.n14251 41.419
R6926 VSS.n14249 VSS.n14247 41.419
R6927 VSS.n17554 VSS.n17552 41.419
R6928 VSS.n17547 VSS.n17544 41.419
R6929 VSS.n17542 VSS.n17539 41.419
R6930 VSS.n17537 VSS.n17535 41.419
R6931 VSS.n17386 VSS.n17384 41.419
R6932 VSS.n17379 VSS.n17376 41.419
R6933 VSS.n17374 VSS.n17371 41.419
R6934 VSS.n17369 VSS.n17367 41.419
R6935 VSS.n17218 VSS.n17216 41.419
R6936 VSS.n17211 VSS.n17208 41.419
R6937 VSS.n17206 VSS.n17203 41.419
R6938 VSS.n17201 VSS.n17199 41.419
R6939 VSS.n17050 VSS.n17048 41.419
R6940 VSS.n17043 VSS.n17040 41.419
R6941 VSS.n17038 VSS.n17035 41.419
R6942 VSS.n17033 VSS.n17031 41.419
R6943 VSS.n16882 VSS.n16880 41.419
R6944 VSS.n16875 VSS.n16872 41.419
R6945 VSS.n16870 VSS.n16867 41.419
R6946 VSS.n16865 VSS.n16863 41.419
R6947 VSS.n16714 VSS.n16712 41.419
R6948 VSS.n16707 VSS.n16704 41.419
R6949 VSS.n16702 VSS.n16699 41.419
R6950 VSS.n16697 VSS.n16695 41.419
R6951 VSS.n14041 VSS.n14039 41.419
R6952 VSS.n14036 VSS.n14033 41.419
R6953 VSS.n14031 VSS.n14028 41.419
R6954 VSS.n14026 VSS.n14024 41.419
R6955 VSS.n13861 VSS.n13859 41.419
R6956 VSS.n13856 VSS.n13853 41.419
R6957 VSS.n13851 VSS.n13848 41.419
R6958 VSS.n13846 VSS.n13844 41.419
R6959 VSS.n13681 VSS.n13679 41.419
R6960 VSS.n13676 VSS.n13673 41.419
R6961 VSS.n13671 VSS.n13668 41.419
R6962 VSS.n13666 VSS.n13664 41.419
R6963 VSS.n13501 VSS.n13499 41.419
R6964 VSS.n13496 VSS.n13493 41.419
R6965 VSS.n13491 VSS.n13488 41.419
R6966 VSS.n13486 VSS.n13484 41.419
R6967 VSS.n13321 VSS.n13319 41.419
R6968 VSS.n13316 VSS.n13313 41.419
R6969 VSS.n13311 VSS.n13308 41.419
R6970 VSS.n13306 VSS.n13304 41.419
R6971 VSS.n13141 VSS.n13139 41.419
R6972 VSS.n13136 VSS.n13133 41.419
R6973 VSS.n13131 VSS.n13128 41.419
R6974 VSS.n13126 VSS.n13124 41.419
R6975 VSS.n12961 VSS.n12959 41.419
R6976 VSS.n12956 VSS.n12953 41.419
R6977 VSS.n12951 VSS.n12948 41.419
R6978 VSS.n12946 VSS.n12944 41.419
R6979 VSS.n12781 VSS.n12779 41.419
R6980 VSS.n12776 VSS.n12773 41.419
R6981 VSS.n12771 VSS.n12768 41.419
R6982 VSS.n12766 VSS.n12764 41.419
R6983 VSS.n9352 VSS.n9350 41.419
R6984 VSS.n9347 VSS.n9344 41.419
R6985 VSS.n9342 VSS.n9339 41.419
R6986 VSS.n9337 VSS.n9335 41.419
R6987 VSS.n9520 VSS.n9518 41.419
R6988 VSS.n9515 VSS.n9512 41.419
R6989 VSS.n9510 VSS.n9507 41.419
R6990 VSS.n9505 VSS.n9503 41.419
R6991 VSS.n9688 VSS.n9686 41.419
R6992 VSS.n9683 VSS.n9680 41.419
R6993 VSS.n9678 VSS.n9675 41.419
R6994 VSS.n9673 VSS.n9671 41.419
R6995 VSS.n9856 VSS.n9854 41.419
R6996 VSS.n9851 VSS.n9848 41.419
R6997 VSS.n9846 VSS.n9843 41.419
R6998 VSS.n9841 VSS.n9839 41.419
R6999 VSS.n10024 VSS.n10022 41.419
R7000 VSS.n10019 VSS.n10016 41.419
R7001 VSS.n10014 VSS.n10011 41.419
R7002 VSS.n10009 VSS.n10007 41.419
R7003 VSS.n10192 VSS.n10190 41.419
R7004 VSS.n10187 VSS.n10184 41.419
R7005 VSS.n10182 VSS.n10179 41.419
R7006 VSS.n10177 VSS.n10175 41.419
R7007 VSS.n10360 VSS.n10358 41.419
R7008 VSS.n10355 VSS.n10352 41.419
R7009 VSS.n10350 VSS.n10347 41.419
R7010 VSS.n10345 VSS.n10343 41.419
R7011 VSS.n10518 VSS.n10516 41.419
R7012 VSS.n10512 VSS.n10509 41.419
R7013 VSS.n10507 VSS.n10504 41.419
R7014 VSS.n10502 VSS.n10500 41.419
R7015 VSS.n2354 VSS.n2299 41.419
R7016 VSS.n2353 VSS.n2297 41.419
R7017 VSS.n2349 VSS.n2296 41.419
R7018 VSS.n2345 VSS.n2295 41.419
R7019 VSS.n2264 VSS.n2209 41.419
R7020 VSS.n2263 VSS.n2207 41.419
R7021 VSS.n2259 VSS.n2206 41.419
R7022 VSS.n2255 VSS.n2205 41.419
R7023 VSS.n2174 VSS.n2119 41.419
R7024 VSS.n2173 VSS.n2117 41.419
R7025 VSS.n2169 VSS.n2116 41.419
R7026 VSS.n2165 VSS.n2115 41.419
R7027 VSS.n2084 VSS.n2029 41.419
R7028 VSS.n2083 VSS.n2027 41.419
R7029 VSS.n2079 VSS.n2026 41.419
R7030 VSS.n2075 VSS.n2025 41.419
R7031 VSS.n1994 VSS.n1939 41.419
R7032 VSS.n1993 VSS.n1937 41.419
R7033 VSS.n1989 VSS.n1936 41.419
R7034 VSS.n1985 VSS.n1935 41.419
R7035 VSS.n1904 VSS.n1849 41.419
R7036 VSS.n1903 VSS.n1847 41.419
R7037 VSS.n1899 VSS.n1846 41.419
R7038 VSS.n1895 VSS.n1845 41.419
R7039 VSS.n1814 VSS.n1759 41.419
R7040 VSS.n1813 VSS.n1757 41.419
R7041 VSS.n1809 VSS.n1756 41.419
R7042 VSS.n1805 VSS.n1755 41.419
R7043 VSS.n1724 VSS.n1669 41.419
R7044 VSS.n1723 VSS.n1667 41.419
R7045 VSS.n1719 VSS.n1666 41.419
R7046 VSS.n1715 VSS.n1665 41.419
R7047 VSS.n6208 VSS.n6090 41.419
R7048 VSS.n6209 VSS.n6088 41.419
R7049 VSS.n6213 VSS.n6087 41.419
R7050 VSS.n6217 VSS.n6086 41.419
R7051 VSS.n6272 VSS.n5974 41.419
R7052 VSS.n6273 VSS.n5972 41.419
R7053 VSS.n6277 VSS.n5971 41.419
R7054 VSS.n6281 VSS.n5970 41.419
R7055 VSS.n6336 VSS.n5858 41.419
R7056 VSS.n6337 VSS.n5856 41.419
R7057 VSS.n6341 VSS.n5855 41.419
R7058 VSS.n6345 VSS.n5854 41.419
R7059 VSS.n6963 VSS.n6962 41.419
R7060 VSS.n6965 VSS.n6964 41.419
R7061 VSS.n6970 VSS.n6969 41.419
R7062 VSS.n6973 VSS.n6972 41.419
R7063 VSS.n6468 VSS.n6413 41.419
R7064 VSS.n6467 VSS.n6411 41.419
R7065 VSS.n6463 VSS.n6410 41.419
R7066 VSS.n6459 VSS.n6409 41.419
R7067 VSS.n6558 VSS.n6503 41.419
R7068 VSS.n6557 VSS.n6501 41.419
R7069 VSS.n6553 VSS.n6500 41.419
R7070 VSS.n6549 VSS.n6499 41.419
R7071 VSS.n6648 VSS.n6593 41.419
R7072 VSS.n6647 VSS.n6591 41.419
R7073 VSS.n6643 VSS.n6590 41.419
R7074 VSS.n6639 VSS.n6589 41.419
R7075 VSS.n17978 VSS.n17932 41.419
R7076 VSS.n17974 VSS.n17933 41.419
R7077 VSS.n17970 VSS.n17934 41.419
R7078 VSS.n17966 VSS.n17935 41.419
R7079 VSS.n14429 VSS.n14428 41.419
R7080 VSS.n14434 VSS.n14433 41.419
R7081 VSS.n14439 VSS.n14438 41.419
R7082 VSS.n14444 VSS.n14443 41.419
R7083 VSS.n14249 VSS.n14248 41.419
R7084 VSS.n14254 VSS.n14253 41.419
R7085 VSS.n14259 VSS.n14258 41.419
R7086 VSS.n14264 VSS.n14263 41.419
R7087 VSS.n17537 VSS.n17536 41.419
R7088 VSS.n17542 VSS.n17541 41.419
R7089 VSS.n17547 VSS.n17546 41.419
R7090 VSS.n17554 VSS.n17553 41.419
R7091 VSS.n17369 VSS.n17368 41.419
R7092 VSS.n17374 VSS.n17373 41.419
R7093 VSS.n17379 VSS.n17378 41.419
R7094 VSS.n17386 VSS.n17385 41.419
R7095 VSS.n17201 VSS.n17200 41.419
R7096 VSS.n17206 VSS.n17205 41.419
R7097 VSS.n17211 VSS.n17210 41.419
R7098 VSS.n17218 VSS.n17217 41.419
R7099 VSS.n17033 VSS.n17032 41.419
R7100 VSS.n17038 VSS.n17037 41.419
R7101 VSS.n17043 VSS.n17042 41.419
R7102 VSS.n17050 VSS.n17049 41.419
R7103 VSS.n16865 VSS.n16864 41.419
R7104 VSS.n16870 VSS.n16869 41.419
R7105 VSS.n16875 VSS.n16874 41.419
R7106 VSS.n16882 VSS.n16881 41.419
R7107 VSS.n16697 VSS.n16696 41.419
R7108 VSS.n16702 VSS.n16701 41.419
R7109 VSS.n16707 VSS.n16706 41.419
R7110 VSS.n16714 VSS.n16713 41.419
R7111 VSS.n14026 VSS.n14025 41.419
R7112 VSS.n14031 VSS.n14030 41.419
R7113 VSS.n14036 VSS.n14035 41.419
R7114 VSS.n14041 VSS.n14040 41.419
R7115 VSS.n13846 VSS.n13845 41.419
R7116 VSS.n13851 VSS.n13850 41.419
R7117 VSS.n13856 VSS.n13855 41.419
R7118 VSS.n13861 VSS.n13860 41.419
R7119 VSS.n13666 VSS.n13665 41.419
R7120 VSS.n13671 VSS.n13670 41.419
R7121 VSS.n13676 VSS.n13675 41.419
R7122 VSS.n13681 VSS.n13680 41.419
R7123 VSS.n13486 VSS.n13485 41.419
R7124 VSS.n13491 VSS.n13490 41.419
R7125 VSS.n13496 VSS.n13495 41.419
R7126 VSS.n13501 VSS.n13500 41.419
R7127 VSS.n13306 VSS.n13305 41.419
R7128 VSS.n13311 VSS.n13310 41.419
R7129 VSS.n13316 VSS.n13315 41.419
R7130 VSS.n13321 VSS.n13320 41.419
R7131 VSS.n13126 VSS.n13125 41.419
R7132 VSS.n13131 VSS.n13130 41.419
R7133 VSS.n13136 VSS.n13135 41.419
R7134 VSS.n13141 VSS.n13140 41.419
R7135 VSS.n12946 VSS.n12945 41.419
R7136 VSS.n12951 VSS.n12950 41.419
R7137 VSS.n12956 VSS.n12955 41.419
R7138 VSS.n12961 VSS.n12960 41.419
R7139 VSS.n12766 VSS.n12765 41.419
R7140 VSS.n12771 VSS.n12770 41.419
R7141 VSS.n12776 VSS.n12775 41.419
R7142 VSS.n12781 VSS.n12780 41.419
R7143 VSS.n9337 VSS.n9336 41.419
R7144 VSS.n9342 VSS.n9341 41.419
R7145 VSS.n9347 VSS.n9346 41.419
R7146 VSS.n9352 VSS.n9351 41.419
R7147 VSS.n9505 VSS.n9504 41.419
R7148 VSS.n9510 VSS.n9509 41.419
R7149 VSS.n9515 VSS.n9514 41.419
R7150 VSS.n9520 VSS.n9519 41.419
R7151 VSS.n9673 VSS.n9672 41.419
R7152 VSS.n9678 VSS.n9677 41.419
R7153 VSS.n9683 VSS.n9682 41.419
R7154 VSS.n9688 VSS.n9687 41.419
R7155 VSS.n9841 VSS.n9840 41.419
R7156 VSS.n9846 VSS.n9845 41.419
R7157 VSS.n9851 VSS.n9850 41.419
R7158 VSS.n9856 VSS.n9855 41.419
R7159 VSS.n10009 VSS.n10008 41.419
R7160 VSS.n10014 VSS.n10013 41.419
R7161 VSS.n10019 VSS.n10018 41.419
R7162 VSS.n10024 VSS.n10023 41.419
R7163 VSS.n10177 VSS.n10176 41.419
R7164 VSS.n10182 VSS.n10181 41.419
R7165 VSS.n10187 VSS.n10186 41.419
R7166 VSS.n10192 VSS.n10191 41.419
R7167 VSS.n10345 VSS.n10344 41.419
R7168 VSS.n10350 VSS.n10349 41.419
R7169 VSS.n10355 VSS.n10354 41.419
R7170 VSS.n10360 VSS.n10359 41.419
R7171 VSS.n10502 VSS.n10501 41.419
R7172 VSS.n10507 VSS.n10506 41.419
R7173 VSS.n10512 VSS.n10511 41.419
R7174 VSS.n10518 VSS.n10517 41.419
R7175 VSS.n2342 VSS.n2295 41.419
R7176 VSS.n2346 VSS.n2296 41.419
R7177 VSS.n2350 VSS.n2297 41.419
R7178 VSS.n2357 VSS.n2299 41.419
R7179 VSS.n2252 VSS.n2205 41.419
R7180 VSS.n2256 VSS.n2206 41.419
R7181 VSS.n2260 VSS.n2207 41.419
R7182 VSS.n2267 VSS.n2209 41.419
R7183 VSS.n2162 VSS.n2115 41.419
R7184 VSS.n2166 VSS.n2116 41.419
R7185 VSS.n2170 VSS.n2117 41.419
R7186 VSS.n2177 VSS.n2119 41.419
R7187 VSS.n2072 VSS.n2025 41.419
R7188 VSS.n2076 VSS.n2026 41.419
R7189 VSS.n2080 VSS.n2027 41.419
R7190 VSS.n2087 VSS.n2029 41.419
R7191 VSS.n1982 VSS.n1935 41.419
R7192 VSS.n1986 VSS.n1936 41.419
R7193 VSS.n1990 VSS.n1937 41.419
R7194 VSS.n1997 VSS.n1939 41.419
R7195 VSS.n1892 VSS.n1845 41.419
R7196 VSS.n1896 VSS.n1846 41.419
R7197 VSS.n1900 VSS.n1847 41.419
R7198 VSS.n1907 VSS.n1849 41.419
R7199 VSS.n1802 VSS.n1755 41.419
R7200 VSS.n1806 VSS.n1756 41.419
R7201 VSS.n1810 VSS.n1757 41.419
R7202 VSS.n1817 VSS.n1759 41.419
R7203 VSS.n1712 VSS.n1665 41.419
R7204 VSS.n1716 VSS.n1666 41.419
R7205 VSS.n1720 VSS.n1667 41.419
R7206 VSS.n1727 VSS.n1669 41.419
R7207 VSS.n6220 VSS.n6086 41.419
R7208 VSS.n6216 VSS.n6087 41.419
R7209 VSS.n6212 VSS.n6088 41.419
R7210 VSS.n6205 VSS.n6090 41.419
R7211 VSS.n6284 VSS.n5970 41.419
R7212 VSS.n6280 VSS.n5971 41.419
R7213 VSS.n6276 VSS.n5972 41.419
R7214 VSS.n6269 VSS.n5974 41.419
R7215 VSS.n6348 VSS.n5854 41.419
R7216 VSS.n6344 VSS.n5855 41.419
R7217 VSS.n6340 VSS.n5856 41.419
R7218 VSS.n6333 VSS.n5858 41.419
R7219 VSS.n6972 VSS.n6390 41.419
R7220 VSS.n6971 VSS.n6970 41.419
R7221 VSS.n6964 VSS.n6392 41.419
R7222 VSS.n6962 VSS.n6961 41.419
R7223 VSS.n6456 VSS.n6409 41.419
R7224 VSS.n6460 VSS.n6410 41.419
R7225 VSS.n6464 VSS.n6411 41.419
R7226 VSS.n6471 VSS.n6413 41.419
R7227 VSS.n6546 VSS.n6499 41.419
R7228 VSS.n6550 VSS.n6500 41.419
R7229 VSS.n6554 VSS.n6501 41.419
R7230 VSS.n6561 VSS.n6503 41.419
R7231 VSS.n6636 VSS.n6589 41.419
R7232 VSS.n6640 VSS.n6590 41.419
R7233 VSS.n6644 VSS.n6591 41.419
R7234 VSS.n6651 VSS.n6593 41.419
R7235 VSS.n17963 VSS.n17935 41.419
R7236 VSS.n17967 VSS.n17934 41.419
R7237 VSS.n17971 VSS.n17933 41.419
R7238 VSS.n17975 VSS.n17932 41.419
R7239 VSS.n14456 VSS.n14455 41.418
R7240 VSS.n14453 VSS.n14452 41.418
R7241 VSS.n14450 VSS.n14449 41.418
R7242 VSS.n14447 VSS.n14446 41.418
R7243 VSS.n14416 VSS.n14414 41.418
R7244 VSS.n14419 VSS.n14417 41.418
R7245 VSS.n14422 VSS.n14420 41.418
R7246 VSS.n14425 VSS.n14423 41.418
R7247 VSS.n14416 VSS.n14415 41.418
R7248 VSS.n14419 VSS.n14418 41.418
R7249 VSS.n14422 VSS.n14421 41.418
R7250 VSS.n14425 VSS.n14424 41.418
R7251 VSS.n14447 VSS.n14445 41.418
R7252 VSS.n14450 VSS.n14448 41.418
R7253 VSS.n14453 VSS.n14451 41.418
R7254 VSS.n14456 VSS.n14454 41.418
R7255 VSS.n14276 VSS.n14275 41.418
R7256 VSS.n14273 VSS.n14272 41.418
R7257 VSS.n14270 VSS.n14269 41.418
R7258 VSS.n14267 VSS.n14266 41.418
R7259 VSS.n14236 VSS.n14234 41.418
R7260 VSS.n14239 VSS.n14237 41.418
R7261 VSS.n14242 VSS.n14240 41.418
R7262 VSS.n14245 VSS.n14243 41.418
R7263 VSS.n14236 VSS.n14235 41.418
R7264 VSS.n14239 VSS.n14238 41.418
R7265 VSS.n14242 VSS.n14241 41.418
R7266 VSS.n14245 VSS.n14244 41.418
R7267 VSS.n14267 VSS.n14265 41.418
R7268 VSS.n14270 VSS.n14268 41.418
R7269 VSS.n14273 VSS.n14271 41.418
R7270 VSS.n14276 VSS.n14274 41.418
R7271 VSS.n17575 VSS.n17574 41.418
R7272 VSS.n17569 VSS.n17568 41.418
R7273 VSS.n17563 VSS.n17562 41.418
R7274 VSS.n17557 VSS.n17556 41.418
R7275 VSS.n17578 VSS.n17576 41.418
R7276 VSS.n17572 VSS.n17570 41.418
R7277 VSS.n17566 VSS.n17564 41.418
R7278 VSS.n17560 VSS.n17558 41.418
R7279 VSS.n17572 VSS.n17571 41.418
R7280 VSS.n17566 VSS.n17565 41.418
R7281 VSS.n17560 VSS.n17559 41.418
R7282 VSS.n17578 VSS.n17577 41.418
R7283 VSS.n17575 VSS.n17573 41.418
R7284 VSS.n17569 VSS.n17567 41.418
R7285 VSS.n17563 VSS.n17561 41.418
R7286 VSS.n17557 VSS.n17555 41.418
R7287 VSS.n17407 VSS.n17406 41.418
R7288 VSS.n17401 VSS.n17400 41.418
R7289 VSS.n17395 VSS.n17394 41.418
R7290 VSS.n17389 VSS.n17388 41.418
R7291 VSS.n17410 VSS.n17408 41.418
R7292 VSS.n17404 VSS.n17402 41.418
R7293 VSS.n17398 VSS.n17396 41.418
R7294 VSS.n17392 VSS.n17390 41.418
R7295 VSS.n17404 VSS.n17403 41.418
R7296 VSS.n17398 VSS.n17397 41.418
R7297 VSS.n17392 VSS.n17391 41.418
R7298 VSS.n17410 VSS.n17409 41.418
R7299 VSS.n17407 VSS.n17405 41.418
R7300 VSS.n17401 VSS.n17399 41.418
R7301 VSS.n17395 VSS.n17393 41.418
R7302 VSS.n17389 VSS.n17387 41.418
R7303 VSS.n17239 VSS.n17238 41.418
R7304 VSS.n17233 VSS.n17232 41.418
R7305 VSS.n17227 VSS.n17226 41.418
R7306 VSS.n17221 VSS.n17220 41.418
R7307 VSS.n17242 VSS.n17240 41.418
R7308 VSS.n17236 VSS.n17234 41.418
R7309 VSS.n17230 VSS.n17228 41.418
R7310 VSS.n17224 VSS.n17222 41.418
R7311 VSS.n17236 VSS.n17235 41.418
R7312 VSS.n17230 VSS.n17229 41.418
R7313 VSS.n17224 VSS.n17223 41.418
R7314 VSS.n17242 VSS.n17241 41.418
R7315 VSS.n17239 VSS.n17237 41.418
R7316 VSS.n17233 VSS.n17231 41.418
R7317 VSS.n17227 VSS.n17225 41.418
R7318 VSS.n17221 VSS.n17219 41.418
R7319 VSS.n17071 VSS.n17070 41.418
R7320 VSS.n17065 VSS.n17064 41.418
R7321 VSS.n17059 VSS.n17058 41.418
R7322 VSS.n17053 VSS.n17052 41.418
R7323 VSS.n17074 VSS.n17072 41.418
R7324 VSS.n17068 VSS.n17066 41.418
R7325 VSS.n17062 VSS.n17060 41.418
R7326 VSS.n17056 VSS.n17054 41.418
R7327 VSS.n17068 VSS.n17067 41.418
R7328 VSS.n17062 VSS.n17061 41.418
R7329 VSS.n17056 VSS.n17055 41.418
R7330 VSS.n17074 VSS.n17073 41.418
R7331 VSS.n17071 VSS.n17069 41.418
R7332 VSS.n17065 VSS.n17063 41.418
R7333 VSS.n17059 VSS.n17057 41.418
R7334 VSS.n17053 VSS.n17051 41.418
R7335 VSS.n16903 VSS.n16902 41.418
R7336 VSS.n16897 VSS.n16896 41.418
R7337 VSS.n16891 VSS.n16890 41.418
R7338 VSS.n16885 VSS.n16884 41.418
R7339 VSS.n16906 VSS.n16904 41.418
R7340 VSS.n16900 VSS.n16898 41.418
R7341 VSS.n16894 VSS.n16892 41.418
R7342 VSS.n16888 VSS.n16886 41.418
R7343 VSS.n16900 VSS.n16899 41.418
R7344 VSS.n16894 VSS.n16893 41.418
R7345 VSS.n16888 VSS.n16887 41.418
R7346 VSS.n16906 VSS.n16905 41.418
R7347 VSS.n16903 VSS.n16901 41.418
R7348 VSS.n16897 VSS.n16895 41.418
R7349 VSS.n16891 VSS.n16889 41.418
R7350 VSS.n16885 VSS.n16883 41.418
R7351 VSS.n16735 VSS.n16734 41.418
R7352 VSS.n16729 VSS.n16728 41.418
R7353 VSS.n16723 VSS.n16722 41.418
R7354 VSS.n16717 VSS.n16716 41.418
R7355 VSS.n16738 VSS.n16736 41.418
R7356 VSS.n16732 VSS.n16730 41.418
R7357 VSS.n16726 VSS.n16724 41.418
R7358 VSS.n16720 VSS.n16718 41.418
R7359 VSS.n16732 VSS.n16731 41.418
R7360 VSS.n16726 VSS.n16725 41.418
R7361 VSS.n16720 VSS.n16719 41.418
R7362 VSS.n16738 VSS.n16737 41.418
R7363 VSS.n16735 VSS.n16733 41.418
R7364 VSS.n16729 VSS.n16727 41.418
R7365 VSS.n16723 VSS.n16721 41.418
R7366 VSS.n16717 VSS.n16715 41.418
R7367 VSS.n14053 VSS.n14052 41.418
R7368 VSS.n14050 VSS.n14049 41.418
R7369 VSS.n14047 VSS.n14046 41.418
R7370 VSS.n14044 VSS.n14043 41.418
R7371 VSS.n14013 VSS.n14011 41.418
R7372 VSS.n14016 VSS.n14014 41.418
R7373 VSS.n14019 VSS.n14017 41.418
R7374 VSS.n14022 VSS.n14020 41.418
R7375 VSS.n14013 VSS.n14012 41.418
R7376 VSS.n14016 VSS.n14015 41.418
R7377 VSS.n14019 VSS.n14018 41.418
R7378 VSS.n14022 VSS.n14021 41.418
R7379 VSS.n14044 VSS.n14042 41.418
R7380 VSS.n14047 VSS.n14045 41.418
R7381 VSS.n14050 VSS.n14048 41.418
R7382 VSS.n14053 VSS.n14051 41.418
R7383 VSS.n13873 VSS.n13872 41.418
R7384 VSS.n13870 VSS.n13869 41.418
R7385 VSS.n13867 VSS.n13866 41.418
R7386 VSS.n13864 VSS.n13863 41.418
R7387 VSS.n13833 VSS.n13831 41.418
R7388 VSS.n13836 VSS.n13834 41.418
R7389 VSS.n13839 VSS.n13837 41.418
R7390 VSS.n13842 VSS.n13840 41.418
R7391 VSS.n13833 VSS.n13832 41.418
R7392 VSS.n13836 VSS.n13835 41.418
R7393 VSS.n13839 VSS.n13838 41.418
R7394 VSS.n13842 VSS.n13841 41.418
R7395 VSS.n13864 VSS.n13862 41.418
R7396 VSS.n13867 VSS.n13865 41.418
R7397 VSS.n13870 VSS.n13868 41.418
R7398 VSS.n13873 VSS.n13871 41.418
R7399 VSS.n13693 VSS.n13692 41.418
R7400 VSS.n13690 VSS.n13689 41.418
R7401 VSS.n13687 VSS.n13686 41.418
R7402 VSS.n13684 VSS.n13683 41.418
R7403 VSS.n13653 VSS.n13651 41.418
R7404 VSS.n13656 VSS.n13654 41.418
R7405 VSS.n13659 VSS.n13657 41.418
R7406 VSS.n13662 VSS.n13660 41.418
R7407 VSS.n13653 VSS.n13652 41.418
R7408 VSS.n13656 VSS.n13655 41.418
R7409 VSS.n13659 VSS.n13658 41.418
R7410 VSS.n13662 VSS.n13661 41.418
R7411 VSS.n13684 VSS.n13682 41.418
R7412 VSS.n13687 VSS.n13685 41.418
R7413 VSS.n13690 VSS.n13688 41.418
R7414 VSS.n13693 VSS.n13691 41.418
R7415 VSS.n13513 VSS.n13512 41.418
R7416 VSS.n13510 VSS.n13509 41.418
R7417 VSS.n13507 VSS.n13506 41.418
R7418 VSS.n13504 VSS.n13503 41.418
R7419 VSS.n13473 VSS.n13471 41.418
R7420 VSS.n13476 VSS.n13474 41.418
R7421 VSS.n13479 VSS.n13477 41.418
R7422 VSS.n13482 VSS.n13480 41.418
R7423 VSS.n13473 VSS.n13472 41.418
R7424 VSS.n13476 VSS.n13475 41.418
R7425 VSS.n13479 VSS.n13478 41.418
R7426 VSS.n13482 VSS.n13481 41.418
R7427 VSS.n13504 VSS.n13502 41.418
R7428 VSS.n13507 VSS.n13505 41.418
R7429 VSS.n13510 VSS.n13508 41.418
R7430 VSS.n13513 VSS.n13511 41.418
R7431 VSS.n13333 VSS.n13332 41.418
R7432 VSS.n13330 VSS.n13329 41.418
R7433 VSS.n13327 VSS.n13326 41.418
R7434 VSS.n13324 VSS.n13323 41.418
R7435 VSS.n13293 VSS.n13291 41.418
R7436 VSS.n13296 VSS.n13294 41.418
R7437 VSS.n13299 VSS.n13297 41.418
R7438 VSS.n13302 VSS.n13300 41.418
R7439 VSS.n13293 VSS.n13292 41.418
R7440 VSS.n13296 VSS.n13295 41.418
R7441 VSS.n13299 VSS.n13298 41.418
R7442 VSS.n13302 VSS.n13301 41.418
R7443 VSS.n13324 VSS.n13322 41.418
R7444 VSS.n13327 VSS.n13325 41.418
R7445 VSS.n13330 VSS.n13328 41.418
R7446 VSS.n13333 VSS.n13331 41.418
R7447 VSS.n13153 VSS.n13152 41.418
R7448 VSS.n13150 VSS.n13149 41.418
R7449 VSS.n13147 VSS.n13146 41.418
R7450 VSS.n13144 VSS.n13143 41.418
R7451 VSS.n13113 VSS.n13111 41.418
R7452 VSS.n13116 VSS.n13114 41.418
R7453 VSS.n13119 VSS.n13117 41.418
R7454 VSS.n13122 VSS.n13120 41.418
R7455 VSS.n13113 VSS.n13112 41.418
R7456 VSS.n13116 VSS.n13115 41.418
R7457 VSS.n13119 VSS.n13118 41.418
R7458 VSS.n13122 VSS.n13121 41.418
R7459 VSS.n13144 VSS.n13142 41.418
R7460 VSS.n13147 VSS.n13145 41.418
R7461 VSS.n13150 VSS.n13148 41.418
R7462 VSS.n13153 VSS.n13151 41.418
R7463 VSS.n12973 VSS.n12972 41.418
R7464 VSS.n12970 VSS.n12969 41.418
R7465 VSS.n12967 VSS.n12966 41.418
R7466 VSS.n12964 VSS.n12963 41.418
R7467 VSS.n12933 VSS.n12931 41.418
R7468 VSS.n12936 VSS.n12934 41.418
R7469 VSS.n12939 VSS.n12937 41.418
R7470 VSS.n12942 VSS.n12940 41.418
R7471 VSS.n12933 VSS.n12932 41.418
R7472 VSS.n12936 VSS.n12935 41.418
R7473 VSS.n12939 VSS.n12938 41.418
R7474 VSS.n12942 VSS.n12941 41.418
R7475 VSS.n12964 VSS.n12962 41.418
R7476 VSS.n12967 VSS.n12965 41.418
R7477 VSS.n12970 VSS.n12968 41.418
R7478 VSS.n12973 VSS.n12971 41.418
R7479 VSS.n12793 VSS.n12792 41.418
R7480 VSS.n12790 VSS.n12789 41.418
R7481 VSS.n12787 VSS.n12786 41.418
R7482 VSS.n12784 VSS.n12783 41.418
R7483 VSS.n12753 VSS.n12751 41.418
R7484 VSS.n12756 VSS.n12754 41.418
R7485 VSS.n12759 VSS.n12757 41.418
R7486 VSS.n12762 VSS.n12760 41.418
R7487 VSS.n12753 VSS.n12752 41.418
R7488 VSS.n12756 VSS.n12755 41.418
R7489 VSS.n12759 VSS.n12758 41.418
R7490 VSS.n12762 VSS.n12761 41.418
R7491 VSS.n12784 VSS.n12782 41.418
R7492 VSS.n12787 VSS.n12785 41.418
R7493 VSS.n12790 VSS.n12788 41.418
R7494 VSS.n12793 VSS.n12791 41.418
R7495 VSS.n9364 VSS.n9363 41.418
R7496 VSS.n9361 VSS.n9360 41.418
R7497 VSS.n9358 VSS.n9357 41.418
R7498 VSS.n9355 VSS.n9354 41.418
R7499 VSS.n9324 VSS.n9322 41.418
R7500 VSS.n9327 VSS.n9325 41.418
R7501 VSS.n9330 VSS.n9328 41.418
R7502 VSS.n9333 VSS.n9331 41.418
R7503 VSS.n9324 VSS.n9323 41.418
R7504 VSS.n9327 VSS.n9326 41.418
R7505 VSS.n9330 VSS.n9329 41.418
R7506 VSS.n9333 VSS.n9332 41.418
R7507 VSS.n9355 VSS.n9353 41.418
R7508 VSS.n9358 VSS.n9356 41.418
R7509 VSS.n9361 VSS.n9359 41.418
R7510 VSS.n9364 VSS.n9362 41.418
R7511 VSS.n9532 VSS.n9531 41.418
R7512 VSS.n9529 VSS.n9528 41.418
R7513 VSS.n9526 VSS.n9525 41.418
R7514 VSS.n9523 VSS.n9522 41.418
R7515 VSS.n9492 VSS.n9490 41.418
R7516 VSS.n9495 VSS.n9493 41.418
R7517 VSS.n9498 VSS.n9496 41.418
R7518 VSS.n9501 VSS.n9499 41.418
R7519 VSS.n9492 VSS.n9491 41.418
R7520 VSS.n9495 VSS.n9494 41.418
R7521 VSS.n9498 VSS.n9497 41.418
R7522 VSS.n9501 VSS.n9500 41.418
R7523 VSS.n9523 VSS.n9521 41.418
R7524 VSS.n9526 VSS.n9524 41.418
R7525 VSS.n9529 VSS.n9527 41.418
R7526 VSS.n9532 VSS.n9530 41.418
R7527 VSS.n9700 VSS.n9699 41.418
R7528 VSS.n9697 VSS.n9696 41.418
R7529 VSS.n9694 VSS.n9693 41.418
R7530 VSS.n9691 VSS.n9690 41.418
R7531 VSS.n9660 VSS.n9658 41.418
R7532 VSS.n9663 VSS.n9661 41.418
R7533 VSS.n9666 VSS.n9664 41.418
R7534 VSS.n9669 VSS.n9667 41.418
R7535 VSS.n9660 VSS.n9659 41.418
R7536 VSS.n9663 VSS.n9662 41.418
R7537 VSS.n9666 VSS.n9665 41.418
R7538 VSS.n9669 VSS.n9668 41.418
R7539 VSS.n9691 VSS.n9689 41.418
R7540 VSS.n9694 VSS.n9692 41.418
R7541 VSS.n9697 VSS.n9695 41.418
R7542 VSS.n9700 VSS.n9698 41.418
R7543 VSS.n9868 VSS.n9867 41.418
R7544 VSS.n9865 VSS.n9864 41.418
R7545 VSS.n9862 VSS.n9861 41.418
R7546 VSS.n9859 VSS.n9858 41.418
R7547 VSS.n9828 VSS.n9826 41.418
R7548 VSS.n9831 VSS.n9829 41.418
R7549 VSS.n9834 VSS.n9832 41.418
R7550 VSS.n9837 VSS.n9835 41.418
R7551 VSS.n9828 VSS.n9827 41.418
R7552 VSS.n9831 VSS.n9830 41.418
R7553 VSS.n9834 VSS.n9833 41.418
R7554 VSS.n9837 VSS.n9836 41.418
R7555 VSS.n9859 VSS.n9857 41.418
R7556 VSS.n9862 VSS.n9860 41.418
R7557 VSS.n9865 VSS.n9863 41.418
R7558 VSS.n9868 VSS.n9866 41.418
R7559 VSS.n10036 VSS.n10035 41.418
R7560 VSS.n10033 VSS.n10032 41.418
R7561 VSS.n10030 VSS.n10029 41.418
R7562 VSS.n10027 VSS.n10026 41.418
R7563 VSS.n9996 VSS.n9994 41.418
R7564 VSS.n9999 VSS.n9997 41.418
R7565 VSS.n10002 VSS.n10000 41.418
R7566 VSS.n10005 VSS.n10003 41.418
R7567 VSS.n9996 VSS.n9995 41.418
R7568 VSS.n9999 VSS.n9998 41.418
R7569 VSS.n10002 VSS.n10001 41.418
R7570 VSS.n10005 VSS.n10004 41.418
R7571 VSS.n10027 VSS.n10025 41.418
R7572 VSS.n10030 VSS.n10028 41.418
R7573 VSS.n10033 VSS.n10031 41.418
R7574 VSS.n10036 VSS.n10034 41.418
R7575 VSS.n10204 VSS.n10203 41.418
R7576 VSS.n10201 VSS.n10200 41.418
R7577 VSS.n10198 VSS.n10197 41.418
R7578 VSS.n10195 VSS.n10194 41.418
R7579 VSS.n10164 VSS.n10162 41.418
R7580 VSS.n10167 VSS.n10165 41.418
R7581 VSS.n10170 VSS.n10168 41.418
R7582 VSS.n10173 VSS.n10171 41.418
R7583 VSS.n10164 VSS.n10163 41.418
R7584 VSS.n10167 VSS.n10166 41.418
R7585 VSS.n10170 VSS.n10169 41.418
R7586 VSS.n10173 VSS.n10172 41.418
R7587 VSS.n10195 VSS.n10193 41.418
R7588 VSS.n10198 VSS.n10196 41.418
R7589 VSS.n10201 VSS.n10199 41.418
R7590 VSS.n10204 VSS.n10202 41.418
R7591 VSS.n10372 VSS.n10371 41.418
R7592 VSS.n10369 VSS.n10368 41.418
R7593 VSS.n10366 VSS.n10365 41.418
R7594 VSS.n10363 VSS.n10362 41.418
R7595 VSS.n10332 VSS.n10330 41.418
R7596 VSS.n10335 VSS.n10333 41.418
R7597 VSS.n10338 VSS.n10336 41.418
R7598 VSS.n10341 VSS.n10339 41.418
R7599 VSS.n10332 VSS.n10331 41.418
R7600 VSS.n10335 VSS.n10334 41.418
R7601 VSS.n10338 VSS.n10337 41.418
R7602 VSS.n10341 VSS.n10340 41.418
R7603 VSS.n10363 VSS.n10361 41.418
R7604 VSS.n10366 VSS.n10364 41.418
R7605 VSS.n10369 VSS.n10367 41.418
R7606 VSS.n10372 VSS.n10370 41.418
R7607 VSS.n10539 VSS.n10538 41.418
R7608 VSS.n10533 VSS.n10532 41.418
R7609 VSS.n10527 VSS.n10526 41.418
R7610 VSS.n10521 VSS.n10520 41.418
R7611 VSS.n10542 VSS.n10540 41.418
R7612 VSS.n10536 VSS.n10534 41.418
R7613 VSS.n10530 VSS.n10528 41.418
R7614 VSS.n10524 VSS.n10522 41.418
R7615 VSS.n10536 VSS.n10535 41.418
R7616 VSS.n10530 VSS.n10529 41.418
R7617 VSS.n10524 VSS.n10523 41.418
R7618 VSS.n10542 VSS.n10541 41.418
R7619 VSS.n10539 VSS.n10537 41.418
R7620 VSS.n10533 VSS.n10531 41.418
R7621 VSS.n10527 VSS.n10525 41.418
R7622 VSS.n10521 VSS.n10519 41.418
R7623 VSS.n2372 VSS.n2303 41.418
R7624 VSS.n2369 VSS.n2302 41.418
R7625 VSS.n2365 VSS.n2301 41.418
R7626 VSS.n2361 VSS.n2300 41.418
R7627 VSS.n2291 VSS.n2289 41.418
R7628 VSS.n2329 VSS.n2292 41.418
R7629 VSS.n2333 VSS.n2293 41.418
R7630 VSS.n2337 VSS.n2294 41.418
R7631 VSS.n2328 VSS.n2291 41.418
R7632 VSS.n2332 VSS.n2292 41.418
R7633 VSS.n2336 VSS.n2293 41.418
R7634 VSS.n2339 VSS.n2294 41.418
R7635 VSS.n2358 VSS.n2300 41.418
R7636 VSS.n2362 VSS.n2301 41.418
R7637 VSS.n2366 VSS.n2302 41.418
R7638 VSS.n2370 VSS.n2303 41.418
R7639 VSS.n2282 VSS.n2213 41.418
R7640 VSS.n2279 VSS.n2212 41.418
R7641 VSS.n2275 VSS.n2211 41.418
R7642 VSS.n2271 VSS.n2210 41.418
R7643 VSS.n2201 VSS.n2199 41.418
R7644 VSS.n2239 VSS.n2202 41.418
R7645 VSS.n2243 VSS.n2203 41.418
R7646 VSS.n2247 VSS.n2204 41.418
R7647 VSS.n2238 VSS.n2201 41.418
R7648 VSS.n2242 VSS.n2202 41.418
R7649 VSS.n2246 VSS.n2203 41.418
R7650 VSS.n2249 VSS.n2204 41.418
R7651 VSS.n2268 VSS.n2210 41.418
R7652 VSS.n2272 VSS.n2211 41.418
R7653 VSS.n2276 VSS.n2212 41.418
R7654 VSS.n2280 VSS.n2213 41.418
R7655 VSS.n2192 VSS.n2123 41.418
R7656 VSS.n2189 VSS.n2122 41.418
R7657 VSS.n2185 VSS.n2121 41.418
R7658 VSS.n2181 VSS.n2120 41.418
R7659 VSS.n2111 VSS.n2109 41.418
R7660 VSS.n2149 VSS.n2112 41.418
R7661 VSS.n2153 VSS.n2113 41.418
R7662 VSS.n2157 VSS.n2114 41.418
R7663 VSS.n2148 VSS.n2111 41.418
R7664 VSS.n2152 VSS.n2112 41.418
R7665 VSS.n2156 VSS.n2113 41.418
R7666 VSS.n2159 VSS.n2114 41.418
R7667 VSS.n2178 VSS.n2120 41.418
R7668 VSS.n2182 VSS.n2121 41.418
R7669 VSS.n2186 VSS.n2122 41.418
R7670 VSS.n2190 VSS.n2123 41.418
R7671 VSS.n2102 VSS.n2033 41.418
R7672 VSS.n2099 VSS.n2032 41.418
R7673 VSS.n2095 VSS.n2031 41.418
R7674 VSS.n2091 VSS.n2030 41.418
R7675 VSS.n2021 VSS.n2019 41.418
R7676 VSS.n2059 VSS.n2022 41.418
R7677 VSS.n2063 VSS.n2023 41.418
R7678 VSS.n2067 VSS.n2024 41.418
R7679 VSS.n2058 VSS.n2021 41.418
R7680 VSS.n2062 VSS.n2022 41.418
R7681 VSS.n2066 VSS.n2023 41.418
R7682 VSS.n2069 VSS.n2024 41.418
R7683 VSS.n2088 VSS.n2030 41.418
R7684 VSS.n2092 VSS.n2031 41.418
R7685 VSS.n2096 VSS.n2032 41.418
R7686 VSS.n2100 VSS.n2033 41.418
R7687 VSS.n2012 VSS.n1943 41.418
R7688 VSS.n2009 VSS.n1942 41.418
R7689 VSS.n2005 VSS.n1941 41.418
R7690 VSS.n2001 VSS.n1940 41.418
R7691 VSS.n1931 VSS.n1929 41.418
R7692 VSS.n1969 VSS.n1932 41.418
R7693 VSS.n1973 VSS.n1933 41.418
R7694 VSS.n1977 VSS.n1934 41.418
R7695 VSS.n1968 VSS.n1931 41.418
R7696 VSS.n1972 VSS.n1932 41.418
R7697 VSS.n1976 VSS.n1933 41.418
R7698 VSS.n1979 VSS.n1934 41.418
R7699 VSS.n1998 VSS.n1940 41.418
R7700 VSS.n2002 VSS.n1941 41.418
R7701 VSS.n2006 VSS.n1942 41.418
R7702 VSS.n2010 VSS.n1943 41.418
R7703 VSS.n1922 VSS.n1853 41.418
R7704 VSS.n1919 VSS.n1852 41.418
R7705 VSS.n1915 VSS.n1851 41.418
R7706 VSS.n1911 VSS.n1850 41.418
R7707 VSS.n1841 VSS.n1839 41.418
R7708 VSS.n1879 VSS.n1842 41.418
R7709 VSS.n1883 VSS.n1843 41.418
R7710 VSS.n1887 VSS.n1844 41.418
R7711 VSS.n1878 VSS.n1841 41.418
R7712 VSS.n1882 VSS.n1842 41.418
R7713 VSS.n1886 VSS.n1843 41.418
R7714 VSS.n1889 VSS.n1844 41.418
R7715 VSS.n1908 VSS.n1850 41.418
R7716 VSS.n1912 VSS.n1851 41.418
R7717 VSS.n1916 VSS.n1852 41.418
R7718 VSS.n1920 VSS.n1853 41.418
R7719 VSS.n1832 VSS.n1763 41.418
R7720 VSS.n1829 VSS.n1762 41.418
R7721 VSS.n1825 VSS.n1761 41.418
R7722 VSS.n1821 VSS.n1760 41.418
R7723 VSS.n1751 VSS.n1749 41.418
R7724 VSS.n1789 VSS.n1752 41.418
R7725 VSS.n1793 VSS.n1753 41.418
R7726 VSS.n1797 VSS.n1754 41.418
R7727 VSS.n1788 VSS.n1751 41.418
R7728 VSS.n1792 VSS.n1752 41.418
R7729 VSS.n1796 VSS.n1753 41.418
R7730 VSS.n1799 VSS.n1754 41.418
R7731 VSS.n1818 VSS.n1760 41.418
R7732 VSS.n1822 VSS.n1761 41.418
R7733 VSS.n1826 VSS.n1762 41.418
R7734 VSS.n1830 VSS.n1763 41.418
R7735 VSS.n1742 VSS.n1673 41.418
R7736 VSS.n1739 VSS.n1672 41.418
R7737 VSS.n1735 VSS.n1671 41.418
R7738 VSS.n1731 VSS.n1670 41.418
R7739 VSS.n1661 VSS.n1659 41.418
R7740 VSS.n1699 VSS.n1662 41.418
R7741 VSS.n1703 VSS.n1663 41.418
R7742 VSS.n1707 VSS.n1664 41.418
R7743 VSS.n1698 VSS.n1661 41.418
R7744 VSS.n1702 VSS.n1662 41.418
R7745 VSS.n1706 VSS.n1663 41.418
R7746 VSS.n1709 VSS.n1664 41.418
R7747 VSS.n1728 VSS.n1670 41.418
R7748 VSS.n1732 VSS.n1671 41.418
R7749 VSS.n1736 VSS.n1672 41.418
R7750 VSS.n1740 VSS.n1673 41.418
R7751 VSS.n6191 VSS.n6097 41.418
R7752 VSS.n6195 VSS.n6095 41.418
R7753 VSS.n6199 VSS.n6093 41.418
R7754 VSS.n6202 VSS.n6091 41.418
R7755 VSS.n6237 VSS.n6098 41.418
R7756 VSS.n6233 VSS.n6096 41.418
R7757 VSS.n6229 VSS.n6094 41.418
R7758 VSS.n6225 VSS.n6092 41.418
R7759 VSS.n6236 VSS.n6096 41.418
R7760 VSS.n6232 VSS.n6094 41.418
R7761 VSS.n6228 VSS.n6092 41.418
R7762 VSS.n6108 VSS.n6098 41.418
R7763 VSS.n6097 VSS.n6076 41.418
R7764 VSS.n6192 VSS.n6095 41.418
R7765 VSS.n6196 VSS.n6093 41.418
R7766 VSS.n6200 VSS.n6091 41.418
R7767 VSS.n6255 VSS.n5981 41.418
R7768 VSS.n6259 VSS.n5979 41.418
R7769 VSS.n6263 VSS.n5977 41.418
R7770 VSS.n6266 VSS.n5975 41.418
R7771 VSS.n6301 VSS.n5982 41.418
R7772 VSS.n6297 VSS.n5980 41.418
R7773 VSS.n6293 VSS.n5978 41.418
R7774 VSS.n6289 VSS.n5976 41.418
R7775 VSS.n6300 VSS.n5980 41.418
R7776 VSS.n6296 VSS.n5978 41.418
R7777 VSS.n6292 VSS.n5976 41.418
R7778 VSS.n5992 VSS.n5982 41.418
R7779 VSS.n5981 VSS.n5960 41.418
R7780 VSS.n6256 VSS.n5979 41.418
R7781 VSS.n6260 VSS.n5977 41.418
R7782 VSS.n6264 VSS.n5975 41.418
R7783 VSS.n6319 VSS.n5865 41.418
R7784 VSS.n6323 VSS.n5863 41.418
R7785 VSS.n6327 VSS.n5861 41.418
R7786 VSS.n6330 VSS.n5859 41.418
R7787 VSS.n6365 VSS.n5866 41.418
R7788 VSS.n6361 VSS.n5864 41.418
R7789 VSS.n6357 VSS.n5862 41.418
R7790 VSS.n6353 VSS.n5860 41.418
R7791 VSS.n6364 VSS.n5864 41.418
R7792 VSS.n6360 VSS.n5862 41.418
R7793 VSS.n6356 VSS.n5860 41.418
R7794 VSS.n5876 VSS.n5866 41.418
R7795 VSS.n5865 VSS.n5844 41.418
R7796 VSS.n6320 VSS.n5863 41.418
R7797 VSS.n6324 VSS.n5861 41.418
R7798 VSS.n6328 VSS.n5859 41.418
R7799 VSS.n6943 VSS.n6398 41.418
R7800 VSS.n6950 VSS.n6949 41.418
R7801 VSS.n6954 VSS.n6396 41.418
R7802 VSS.n6957 VSS.n6956 41.418
R7803 VSS.n6992 VSS.n6991 41.418
R7804 VSS.n6987 VSS.n6386 41.418
R7805 VSS.n6985 VSS.n6984 41.418
R7806 VSS.n6980 VSS.n6389 41.418
R7807 VSS.n6386 VSS.n6384 41.418
R7808 VSS.n6986 VSS.n6985 41.418
R7809 VSS.n6389 VSS.n6387 41.418
R7810 VSS.n6993 VSS.n6992 41.418
R7811 VSS.n6944 VSS.n6943 41.418
R7812 VSS.n6949 VSS.n6948 41.418
R7813 VSS.n6951 VSS.n6396 41.418
R7814 VSS.n6956 VSS.n6955 41.418
R7815 VSS.n6486 VSS.n6417 41.418
R7816 VSS.n6483 VSS.n6416 41.418
R7817 VSS.n6479 VSS.n6415 41.418
R7818 VSS.n6475 VSS.n6414 41.418
R7819 VSS.n6405 VSS.n6403 41.418
R7820 VSS.n6443 VSS.n6406 41.418
R7821 VSS.n6447 VSS.n6407 41.418
R7822 VSS.n6451 VSS.n6408 41.418
R7823 VSS.n6442 VSS.n6405 41.418
R7824 VSS.n6446 VSS.n6406 41.418
R7825 VSS.n6450 VSS.n6407 41.418
R7826 VSS.n6453 VSS.n6408 41.418
R7827 VSS.n6472 VSS.n6414 41.418
R7828 VSS.n6476 VSS.n6415 41.418
R7829 VSS.n6480 VSS.n6416 41.418
R7830 VSS.n6484 VSS.n6417 41.418
R7831 VSS.n6576 VSS.n6507 41.418
R7832 VSS.n6573 VSS.n6506 41.418
R7833 VSS.n6569 VSS.n6505 41.418
R7834 VSS.n6565 VSS.n6504 41.418
R7835 VSS.n6495 VSS.n6493 41.418
R7836 VSS.n6533 VSS.n6496 41.418
R7837 VSS.n6537 VSS.n6497 41.418
R7838 VSS.n6541 VSS.n6498 41.418
R7839 VSS.n6532 VSS.n6495 41.418
R7840 VSS.n6536 VSS.n6496 41.418
R7841 VSS.n6540 VSS.n6497 41.418
R7842 VSS.n6543 VSS.n6498 41.418
R7843 VSS.n6562 VSS.n6504 41.418
R7844 VSS.n6566 VSS.n6505 41.418
R7845 VSS.n6570 VSS.n6506 41.418
R7846 VSS.n6574 VSS.n6507 41.418
R7847 VSS.n6666 VSS.n6597 41.418
R7848 VSS.n6663 VSS.n6596 41.418
R7849 VSS.n6659 VSS.n6595 41.418
R7850 VSS.n6655 VSS.n6594 41.418
R7851 VSS.n6585 VSS.n6583 41.418
R7852 VSS.n6623 VSS.n6586 41.418
R7853 VSS.n6627 VSS.n6587 41.418
R7854 VSS.n6631 VSS.n6588 41.418
R7855 VSS.n6622 VSS.n6585 41.418
R7856 VSS.n6626 VSS.n6586 41.418
R7857 VSS.n6630 VSS.n6587 41.418
R7858 VSS.n6633 VSS.n6588 41.418
R7859 VSS.n6652 VSS.n6594 41.418
R7860 VSS.n6656 VSS.n6595 41.418
R7861 VSS.n6660 VSS.n6596 41.418
R7862 VSS.n6664 VSS.n6597 41.418
R7863 VSS.n17991 VSS.n17937 41.418
R7864 VSS.n17990 VSS.n17926 41.418
R7865 VSS.n17986 VSS.n17928 41.418
R7866 VSS.n17982 VSS.n17930 41.418
R7867 VSS.n17954 VSS.n17929 41.418
R7868 VSS.n17958 VSS.n17931 41.418
R7869 VSS.n17994 VSS.n17937 41.418
R7870 VSS.n17987 VSS.n17926 41.418
R7871 VSS.n17983 VSS.n17928 41.418
R7872 VSS.n17979 VSS.n17930 41.418
R7873 VSS.n17951 VSS.n17929 41.418
R7874 VSS.n17955 VSS.n17931 41.418
R7875 VSS.t78 VSS.n17945 40.03
R7876 VSS.t78 VSS.n17938 38.819
R7877 VSS.n17995 VSS.n17938 34.273
R7878 VSS VSS.n342 33.172
R7879 VSS VSS.n18293 33.099
R7880 VSS.n18011 VSS.n17945 32.457
R7881 VSS.n405 VSS.n404 31.034
R7882 VSS.n406 VSS.n357 31.034
R7883 VSS.n18197 VSS.n18196 31.034
R7884 VSS.n18198 VSS.n18149 31.034
R7885 VSS.n17950 VSS.n17927 28.99
R7886 VSS.n14468 VSS.n14467 27.554
R7887 VSS.n14288 VSS.n14287 27.554
R7888 VSS.n14482 VSS.n14481 27.554
R7889 VSS.n14494 VSS.n14493 27.554
R7890 VSS.n14506 VSS.n14505 27.554
R7891 VSS.n14518 VSS.n14517 27.554
R7892 VSS.n14530 VSS.n14529 27.554
R7893 VSS.n14542 VSS.n14541 27.554
R7894 VSS.n14066 VSS.n14065 27.554
R7895 VSS.n13885 VSS.n13884 27.554
R7896 VSS.n13705 VSS.n13704 27.554
R7897 VSS.n13525 VSS.n13524 27.554
R7898 VSS.n13345 VSS.n13344 27.554
R7899 VSS.n13165 VSS.n13164 27.554
R7900 VSS.n12985 VSS.n12984 27.554
R7901 VSS.n12805 VSS.n12804 27.554
R7902 VSS.n9209 VSS.n9208 27.554
R7903 VSS.n9377 VSS.n9376 27.554
R7904 VSS.n9545 VSS.n9544 27.554
R7905 VSS.n9713 VSS.n9712 27.554
R7906 VSS.n9881 VSS.n9880 27.554
R7907 VSS.n10049 VSS.n10048 27.554
R7908 VSS.n10217 VSS.n10216 27.554
R7909 VSS.n10385 VSS.n10384 27.554
R7910 VSS.n2341 VSS.n2340 27.554
R7911 VSS.n2251 VSS.n2250 27.554
R7912 VSS.n2161 VSS.n2160 27.554
R7913 VSS.n2071 VSS.n2070 27.554
R7914 VSS.n1981 VSS.n1980 27.554
R7915 VSS.n1891 VSS.n1890 27.554
R7916 VSS.n1801 VSS.n1800 27.554
R7917 VSS.n1711 VSS.n1710 27.554
R7918 VSS.n6223 VSS.n6222 27.554
R7919 VSS.n6287 VSS.n6286 27.554
R7920 VSS.n6351 VSS.n6350 27.554
R7921 VSS.n6976 VSS.n6388 27.554
R7922 VSS.n6455 VSS.n6454 27.554
R7923 VSS.n6545 VSS.n6544 27.554
R7924 VSS.n6635 VSS.n6634 27.554
R7925 VSS.n17961 VSS.n17960 27.554
R7926 VSS.n18090 VSS 27.3
R7927 VSS.n395 VSS.n394 26.896
R7928 VSS.n413 VSS.n353 26.896
R7929 VSS.n18187 VSS.n18186 26.896
R7930 VSS.n18205 VSS.n18143 26.896
R7931 VSS.n14301 VSS.n14300 26.666
R7932 VSS.n14122 VSS.n14121 26.666
R7933 VSS.n17587 VSS.n17586 26.666
R7934 VSS.n17419 VSS.n17418 26.666
R7935 VSS.n17251 VSS.n17250 26.666
R7936 VSS.n17083 VSS.n17082 26.666
R7937 VSS.n16915 VSS.n16914 26.666
R7938 VSS.n16747 VSS.n16746 26.666
R7939 VSS.n13898 VSS.n13897 26.666
R7940 VSS.n13718 VSS.n13717 26.666
R7941 VSS.n13538 VSS.n13537 26.666
R7942 VSS.n13358 VSS.n13357 26.666
R7943 VSS.n13178 VSS.n13177 26.666
R7944 VSS.n12998 VSS.n12997 26.666
R7945 VSS.n12818 VSS.n12817 26.666
R7946 VSS.n12639 VSS.n12638 26.666
R7947 VSS.n7158 VSS.n7157 26.666
R7948 VSS.n7146 VSS.n7145 26.666
R7949 VSS.n7134 VSS.n7133 26.666
R7950 VSS.n7122 VSS.n7121 26.666
R7951 VSS.n7110 VSS.n7109 26.666
R7952 VSS.n7098 VSS.n7097 26.666
R7953 VSS.n7086 VSS.n7085 26.666
R7954 VSS.n10553 VSS.n10552 26.666
R7955 VSS.n2359 VSS.n2356 26.666
R7956 VSS.n2269 VSS.n2266 26.666
R7957 VSS.n2179 VSS.n2176 26.666
R7958 VSS.n2089 VSS.n2086 26.666
R7959 VSS.n1999 VSS.n1996 26.666
R7960 VSS.n1909 VSS.n1906 26.666
R7961 VSS.n1819 VSS.n1816 26.666
R7962 VSS.n1729 VSS.n1726 26.666
R7963 VSS.n6206 VSS.n6204 26.666
R7964 VSS.n6270 VSS.n6268 26.666
R7965 VSS.n6334 VSS.n6332 26.666
R7966 VSS.n6960 VSS.n6959 26.666
R7967 VSS.n6473 VSS.n6470 26.666
R7968 VSS.n6563 VSS.n6560 26.666
R7969 VSS.n6653 VSS.n6650 26.666
R7970 VSS.n18014 VSS.n18013 26.666
R7971 VSS.t10 VSS.n14439 25.542
R7972 VSS.t10 VSS.n14434 25.542
R7973 VSS.t10 VSS.n14429 25.542
R7974 VSS.t10 VSS.n14444 25.542
R7975 VSS.t8 VSS.n14259 25.542
R7976 VSS.t8 VSS.n14254 25.542
R7977 VSS.t8 VSS.n14249 25.542
R7978 VSS.t8 VSS.n14264 25.542
R7979 VSS.t6 VSS.n17547 25.542
R7980 VSS.t6 VSS.n17542 25.542
R7981 VSS.t6 VSS.n17537 25.542
R7982 VSS.t6 VSS.n17554 25.542
R7983 VSS.t2 VSS.n17379 25.542
R7984 VSS.t2 VSS.n17374 25.542
R7985 VSS.t2 VSS.n17369 25.542
R7986 VSS.t2 VSS.n17386 25.542
R7987 VSS.t4 VSS.n17211 25.542
R7988 VSS.t4 VSS.n17206 25.542
R7989 VSS.t4 VSS.n17201 25.542
R7990 VSS.t4 VSS.n17218 25.542
R7991 VSS.t12 VSS.n17043 25.542
R7992 VSS.t12 VSS.n17038 25.542
R7993 VSS.t12 VSS.n17033 25.542
R7994 VSS.t12 VSS.n17050 25.542
R7995 VSS.t14 VSS.n16875 25.542
R7996 VSS.t14 VSS.n16870 25.542
R7997 VSS.t14 VSS.n16865 25.542
R7998 VSS.t14 VSS.n16882 25.542
R7999 VSS.t0 VSS.n16707 25.542
R8000 VSS.t0 VSS.n16702 25.542
R8001 VSS.t0 VSS.n16697 25.542
R8002 VSS.t0 VSS.n16714 25.542
R8003 VSS.t32 VSS.n14036 25.542
R8004 VSS.t32 VSS.n14031 25.542
R8005 VSS.t32 VSS.n14026 25.542
R8006 VSS.t32 VSS.n14041 25.542
R8007 VSS.t46 VSS.n13856 25.542
R8008 VSS.t46 VSS.n13851 25.542
R8009 VSS.t46 VSS.n13846 25.542
R8010 VSS.t46 VSS.n13861 25.542
R8011 VSS.t44 VSS.n13676 25.542
R8012 VSS.t44 VSS.n13671 25.542
R8013 VSS.t44 VSS.n13666 25.542
R8014 VSS.t44 VSS.n13681 25.542
R8015 VSS.t36 VSS.n13496 25.542
R8016 VSS.t36 VSS.n13491 25.542
R8017 VSS.t36 VSS.n13486 25.542
R8018 VSS.t36 VSS.n13501 25.542
R8019 VSS.t34 VSS.n13316 25.542
R8020 VSS.t34 VSS.n13311 25.542
R8021 VSS.t34 VSS.n13306 25.542
R8022 VSS.t34 VSS.n13321 25.542
R8023 VSS.t38 VSS.n13136 25.542
R8024 VSS.t38 VSS.n13131 25.542
R8025 VSS.t38 VSS.n13126 25.542
R8026 VSS.t38 VSS.n13141 25.542
R8027 VSS.t42 VSS.n12956 25.542
R8028 VSS.t42 VSS.n12951 25.542
R8029 VSS.t42 VSS.n12946 25.542
R8030 VSS.t42 VSS.n12961 25.542
R8031 VSS.t40 VSS.n12776 25.542
R8032 VSS.t40 VSS.n12771 25.542
R8033 VSS.t40 VSS.n12766 25.542
R8034 VSS.t40 VSS.n12781 25.542
R8035 VSS.t48 VSS.n9347 25.542
R8036 VSS.t48 VSS.n9342 25.542
R8037 VSS.t48 VSS.n9337 25.542
R8038 VSS.t48 VSS.n9352 25.542
R8039 VSS.t62 VSS.n9515 25.542
R8040 VSS.t62 VSS.n9510 25.542
R8041 VSS.t62 VSS.n9505 25.542
R8042 VSS.t62 VSS.n9520 25.542
R8043 VSS.t60 VSS.n9683 25.542
R8044 VSS.t60 VSS.n9678 25.542
R8045 VSS.t60 VSS.n9673 25.542
R8046 VSS.t60 VSS.n9688 25.542
R8047 VSS.t52 VSS.n9851 25.542
R8048 VSS.t52 VSS.n9846 25.542
R8049 VSS.t52 VSS.n9841 25.542
R8050 VSS.t52 VSS.n9856 25.542
R8051 VSS.t50 VSS.n10019 25.542
R8052 VSS.t50 VSS.n10014 25.542
R8053 VSS.t50 VSS.n10009 25.542
R8054 VSS.t50 VSS.n10024 25.542
R8055 VSS.t54 VSS.n10187 25.542
R8056 VSS.t54 VSS.n10182 25.542
R8057 VSS.t54 VSS.n10177 25.542
R8058 VSS.t54 VSS.n10192 25.542
R8059 VSS.t58 VSS.n10355 25.542
R8060 VSS.t58 VSS.n10350 25.542
R8061 VSS.t58 VSS.n10345 25.542
R8062 VSS.t58 VSS.n10360 25.542
R8063 VSS.t56 VSS.n10512 25.542
R8064 VSS.t56 VSS.n10507 25.542
R8065 VSS.t56 VSS.n10502 25.542
R8066 VSS.t56 VSS.n10518 25.542
R8067 VSS.t24 VSS.n2297 25.542
R8068 VSS.t24 VSS.n2296 25.542
R8069 VSS.t24 VSS.n2295 25.542
R8070 VSS.t24 VSS.n2299 25.542
R8071 VSS.t26 VSS.n2207 25.542
R8072 VSS.t26 VSS.n2206 25.542
R8073 VSS.t26 VSS.n2205 25.542
R8074 VSS.t26 VSS.n2209 25.542
R8075 VSS.t22 VSS.n2117 25.542
R8076 VSS.t22 VSS.n2116 25.542
R8077 VSS.t22 VSS.n2115 25.542
R8078 VSS.t22 VSS.n2119 25.542
R8079 VSS.t18 VSS.n2027 25.542
R8080 VSS.t18 VSS.n2026 25.542
R8081 VSS.t18 VSS.n2025 25.542
R8082 VSS.t18 VSS.n2029 25.542
R8083 VSS.t20 VSS.n1937 25.542
R8084 VSS.t20 VSS.n1936 25.542
R8085 VSS.t20 VSS.n1935 25.542
R8086 VSS.t20 VSS.n1939 25.542
R8087 VSS.t28 VSS.n1847 25.542
R8088 VSS.t28 VSS.n1846 25.542
R8089 VSS.t28 VSS.n1845 25.542
R8090 VSS.t28 VSS.n1849 25.542
R8091 VSS.t30 VSS.n1757 25.542
R8092 VSS.t30 VSS.n1756 25.542
R8093 VSS.t30 VSS.n1755 25.542
R8094 VSS.t30 VSS.n1759 25.542
R8095 VSS.t16 VSS.n1667 25.542
R8096 VSS.t16 VSS.n1666 25.542
R8097 VSS.t16 VSS.n1665 25.542
R8098 VSS.t16 VSS.n1669 25.542
R8099 VSS.t64 VSS.n6088 25.542
R8100 VSS.t64 VSS.n6087 25.542
R8101 VSS.t64 VSS.n6086 25.542
R8102 VSS.t64 VSS.n6090 25.542
R8103 VSS.t76 VSS.n5972 25.542
R8104 VSS.t76 VSS.n5971 25.542
R8105 VSS.t76 VSS.n5970 25.542
R8106 VSS.t76 VSS.n5974 25.542
R8107 VSS.t74 VSS.n5856 25.542
R8108 VSS.t74 VSS.n5855 25.542
R8109 VSS.t74 VSS.n5854 25.542
R8110 VSS.t74 VSS.n5858 25.542
R8111 VSS.n6964 VSS.t68 25.542
R8112 VSS.n6970 VSS.t68 25.542
R8113 VSS.n6972 VSS.t68 25.542
R8114 VSS.n6962 VSS.t68 25.542
R8115 VSS.t66 VSS.n6411 25.542
R8116 VSS.t66 VSS.n6410 25.542
R8117 VSS.t66 VSS.n6409 25.542
R8118 VSS.t66 VSS.n6413 25.542
R8119 VSS.t70 VSS.n6501 25.542
R8120 VSS.t70 VSS.n6500 25.542
R8121 VSS.t70 VSS.n6499 25.542
R8122 VSS.t70 VSS.n6503 25.542
R8123 VSS.t72 VSS.n6591 25.542
R8124 VSS.t72 VSS.n6590 25.542
R8125 VSS.t72 VSS.n6589 25.542
R8126 VSS.t72 VSS.n6593 25.542
R8127 VSS.t78 VSS.n17932 25.542
R8128 VSS.t78 VSS.n17933 25.542
R8129 VSS.t78 VSS.n17934 25.542
R8130 VSS.t78 VSS.n17935 25.542
R8131 VSS.t10 VSS.n14416 25.542
R8132 VSS.t10 VSS.n14419 25.542
R8133 VSS.t10 VSS.n14422 25.542
R8134 VSS.t10 VSS.n14425 25.542
R8135 VSS.t10 VSS.n14447 25.542
R8136 VSS.t10 VSS.n14450 25.542
R8137 VSS.t10 VSS.n14453 25.542
R8138 VSS.t10 VSS.n14456 25.542
R8139 VSS.t8 VSS.n14236 25.542
R8140 VSS.t8 VSS.n14239 25.542
R8141 VSS.t8 VSS.n14242 25.542
R8142 VSS.t8 VSS.n14245 25.542
R8143 VSS.t8 VSS.n14267 25.542
R8144 VSS.t8 VSS.n14270 25.542
R8145 VSS.t8 VSS.n14273 25.542
R8146 VSS.t8 VSS.n14276 25.542
R8147 VSS.t6 VSS.n17578 25.542
R8148 VSS.t6 VSS.n17572 25.542
R8149 VSS.t6 VSS.n17566 25.542
R8150 VSS.t6 VSS.n17560 25.542
R8151 VSS.t6 VSS.n17575 25.542
R8152 VSS.t6 VSS.n17569 25.542
R8153 VSS.t6 VSS.n17563 25.542
R8154 VSS.t6 VSS.n17557 25.542
R8155 VSS.t2 VSS.n17410 25.542
R8156 VSS.t2 VSS.n17404 25.542
R8157 VSS.t2 VSS.n17398 25.542
R8158 VSS.t2 VSS.n17392 25.542
R8159 VSS.t2 VSS.n17407 25.542
R8160 VSS.t2 VSS.n17401 25.542
R8161 VSS.t2 VSS.n17395 25.542
R8162 VSS.t2 VSS.n17389 25.542
R8163 VSS.t4 VSS.n17242 25.542
R8164 VSS.t4 VSS.n17236 25.542
R8165 VSS.t4 VSS.n17230 25.542
R8166 VSS.t4 VSS.n17224 25.542
R8167 VSS.t4 VSS.n17239 25.542
R8168 VSS.t4 VSS.n17233 25.542
R8169 VSS.t4 VSS.n17227 25.542
R8170 VSS.t4 VSS.n17221 25.542
R8171 VSS.t12 VSS.n17074 25.542
R8172 VSS.t12 VSS.n17068 25.542
R8173 VSS.t12 VSS.n17062 25.542
R8174 VSS.t12 VSS.n17056 25.542
R8175 VSS.t12 VSS.n17071 25.542
R8176 VSS.t12 VSS.n17065 25.542
R8177 VSS.t12 VSS.n17059 25.542
R8178 VSS.t12 VSS.n17053 25.542
R8179 VSS.t14 VSS.n16906 25.542
R8180 VSS.t14 VSS.n16900 25.542
R8181 VSS.t14 VSS.n16894 25.542
R8182 VSS.t14 VSS.n16888 25.542
R8183 VSS.t14 VSS.n16903 25.542
R8184 VSS.t14 VSS.n16897 25.542
R8185 VSS.t14 VSS.n16891 25.542
R8186 VSS.t14 VSS.n16885 25.542
R8187 VSS.t0 VSS.n16738 25.542
R8188 VSS.t0 VSS.n16732 25.542
R8189 VSS.t0 VSS.n16726 25.542
R8190 VSS.t0 VSS.n16720 25.542
R8191 VSS.t0 VSS.n16735 25.542
R8192 VSS.t0 VSS.n16729 25.542
R8193 VSS.t0 VSS.n16723 25.542
R8194 VSS.t0 VSS.n16717 25.542
R8195 VSS.t32 VSS.n14013 25.542
R8196 VSS.t32 VSS.n14016 25.542
R8197 VSS.t32 VSS.n14019 25.542
R8198 VSS.t32 VSS.n14022 25.542
R8199 VSS.t32 VSS.n14044 25.542
R8200 VSS.t32 VSS.n14047 25.542
R8201 VSS.t32 VSS.n14050 25.542
R8202 VSS.t32 VSS.n14053 25.542
R8203 VSS.t46 VSS.n13833 25.542
R8204 VSS.t46 VSS.n13836 25.542
R8205 VSS.t46 VSS.n13839 25.542
R8206 VSS.t46 VSS.n13842 25.542
R8207 VSS.t46 VSS.n13864 25.542
R8208 VSS.t46 VSS.n13867 25.542
R8209 VSS.t46 VSS.n13870 25.542
R8210 VSS.t46 VSS.n13873 25.542
R8211 VSS.t44 VSS.n13653 25.542
R8212 VSS.t44 VSS.n13656 25.542
R8213 VSS.t44 VSS.n13659 25.542
R8214 VSS.t44 VSS.n13662 25.542
R8215 VSS.t44 VSS.n13684 25.542
R8216 VSS.t44 VSS.n13687 25.542
R8217 VSS.t44 VSS.n13690 25.542
R8218 VSS.t44 VSS.n13693 25.542
R8219 VSS.t36 VSS.n13473 25.542
R8220 VSS.t36 VSS.n13476 25.542
R8221 VSS.t36 VSS.n13479 25.542
R8222 VSS.t36 VSS.n13482 25.542
R8223 VSS.t36 VSS.n13504 25.542
R8224 VSS.t36 VSS.n13507 25.542
R8225 VSS.t36 VSS.n13510 25.542
R8226 VSS.t36 VSS.n13513 25.542
R8227 VSS.t34 VSS.n13293 25.542
R8228 VSS.t34 VSS.n13296 25.542
R8229 VSS.t34 VSS.n13299 25.542
R8230 VSS.t34 VSS.n13302 25.542
R8231 VSS.t34 VSS.n13324 25.542
R8232 VSS.t34 VSS.n13327 25.542
R8233 VSS.t34 VSS.n13330 25.542
R8234 VSS.t34 VSS.n13333 25.542
R8235 VSS.t38 VSS.n13113 25.542
R8236 VSS.t38 VSS.n13116 25.542
R8237 VSS.t38 VSS.n13119 25.542
R8238 VSS.t38 VSS.n13122 25.542
R8239 VSS.t38 VSS.n13144 25.542
R8240 VSS.t38 VSS.n13147 25.542
R8241 VSS.t38 VSS.n13150 25.542
R8242 VSS.t38 VSS.n13153 25.542
R8243 VSS.t42 VSS.n12933 25.542
R8244 VSS.t42 VSS.n12936 25.542
R8245 VSS.t42 VSS.n12939 25.542
R8246 VSS.t42 VSS.n12942 25.542
R8247 VSS.t42 VSS.n12964 25.542
R8248 VSS.t42 VSS.n12967 25.542
R8249 VSS.t42 VSS.n12970 25.542
R8250 VSS.t42 VSS.n12973 25.542
R8251 VSS.t40 VSS.n12753 25.542
R8252 VSS.t40 VSS.n12756 25.542
R8253 VSS.t40 VSS.n12759 25.542
R8254 VSS.t40 VSS.n12762 25.542
R8255 VSS.t40 VSS.n12784 25.542
R8256 VSS.t40 VSS.n12787 25.542
R8257 VSS.t40 VSS.n12790 25.542
R8258 VSS.t40 VSS.n12793 25.542
R8259 VSS.t48 VSS.n9324 25.542
R8260 VSS.t48 VSS.n9327 25.542
R8261 VSS.t48 VSS.n9330 25.542
R8262 VSS.t48 VSS.n9333 25.542
R8263 VSS.t48 VSS.n9355 25.542
R8264 VSS.t48 VSS.n9358 25.542
R8265 VSS.t48 VSS.n9361 25.542
R8266 VSS.t48 VSS.n9364 25.542
R8267 VSS.t62 VSS.n9492 25.542
R8268 VSS.t62 VSS.n9495 25.542
R8269 VSS.t62 VSS.n9498 25.542
R8270 VSS.t62 VSS.n9501 25.542
R8271 VSS.t62 VSS.n9523 25.542
R8272 VSS.t62 VSS.n9526 25.542
R8273 VSS.t62 VSS.n9529 25.542
R8274 VSS.t62 VSS.n9532 25.542
R8275 VSS.t60 VSS.n9660 25.542
R8276 VSS.t60 VSS.n9663 25.542
R8277 VSS.t60 VSS.n9666 25.542
R8278 VSS.t60 VSS.n9669 25.542
R8279 VSS.t60 VSS.n9691 25.542
R8280 VSS.t60 VSS.n9694 25.542
R8281 VSS.t60 VSS.n9697 25.542
R8282 VSS.t60 VSS.n9700 25.542
R8283 VSS.t52 VSS.n9828 25.542
R8284 VSS.t52 VSS.n9831 25.542
R8285 VSS.t52 VSS.n9834 25.542
R8286 VSS.t52 VSS.n9837 25.542
R8287 VSS.t52 VSS.n9859 25.542
R8288 VSS.t52 VSS.n9862 25.542
R8289 VSS.t52 VSS.n9865 25.542
R8290 VSS.t52 VSS.n9868 25.542
R8291 VSS.t50 VSS.n9996 25.542
R8292 VSS.t50 VSS.n9999 25.542
R8293 VSS.t50 VSS.n10002 25.542
R8294 VSS.t50 VSS.n10005 25.542
R8295 VSS.t50 VSS.n10027 25.542
R8296 VSS.t50 VSS.n10030 25.542
R8297 VSS.t50 VSS.n10033 25.542
R8298 VSS.t50 VSS.n10036 25.542
R8299 VSS.t54 VSS.n10164 25.542
R8300 VSS.t54 VSS.n10167 25.542
R8301 VSS.t54 VSS.n10170 25.542
R8302 VSS.t54 VSS.n10173 25.542
R8303 VSS.t54 VSS.n10195 25.542
R8304 VSS.t54 VSS.n10198 25.542
R8305 VSS.t54 VSS.n10201 25.542
R8306 VSS.t54 VSS.n10204 25.542
R8307 VSS.t58 VSS.n10332 25.542
R8308 VSS.t58 VSS.n10335 25.542
R8309 VSS.t58 VSS.n10338 25.542
R8310 VSS.t58 VSS.n10341 25.542
R8311 VSS.t58 VSS.n10363 25.542
R8312 VSS.t58 VSS.n10366 25.542
R8313 VSS.t58 VSS.n10369 25.542
R8314 VSS.t58 VSS.n10372 25.542
R8315 VSS.t56 VSS.n10542 25.542
R8316 VSS.t56 VSS.n10536 25.542
R8317 VSS.t56 VSS.n10530 25.542
R8318 VSS.t56 VSS.n10524 25.542
R8319 VSS.t56 VSS.n10539 25.542
R8320 VSS.t56 VSS.n10533 25.542
R8321 VSS.t56 VSS.n10527 25.542
R8322 VSS.t56 VSS.n10521 25.542
R8323 VSS.t24 VSS.n2291 25.542
R8324 VSS.t24 VSS.n2292 25.542
R8325 VSS.t24 VSS.n2293 25.542
R8326 VSS.t24 VSS.n2294 25.542
R8327 VSS.t24 VSS.n2300 25.542
R8328 VSS.t24 VSS.n2301 25.542
R8329 VSS.t24 VSS.n2302 25.542
R8330 VSS.t24 VSS.n2303 25.542
R8331 VSS.t26 VSS.n2201 25.542
R8332 VSS.t26 VSS.n2202 25.542
R8333 VSS.t26 VSS.n2203 25.542
R8334 VSS.t26 VSS.n2204 25.542
R8335 VSS.t26 VSS.n2210 25.542
R8336 VSS.t26 VSS.n2211 25.542
R8337 VSS.t26 VSS.n2212 25.542
R8338 VSS.t26 VSS.n2213 25.542
R8339 VSS.t22 VSS.n2111 25.542
R8340 VSS.t22 VSS.n2112 25.542
R8341 VSS.t22 VSS.n2113 25.542
R8342 VSS.t22 VSS.n2114 25.542
R8343 VSS.t22 VSS.n2120 25.542
R8344 VSS.t22 VSS.n2121 25.542
R8345 VSS.t22 VSS.n2122 25.542
R8346 VSS.t22 VSS.n2123 25.542
R8347 VSS.t18 VSS.n2021 25.542
R8348 VSS.t18 VSS.n2022 25.542
R8349 VSS.t18 VSS.n2023 25.542
R8350 VSS.t18 VSS.n2024 25.542
R8351 VSS.t18 VSS.n2030 25.542
R8352 VSS.t18 VSS.n2031 25.542
R8353 VSS.t18 VSS.n2032 25.542
R8354 VSS.t18 VSS.n2033 25.542
R8355 VSS.t20 VSS.n1931 25.542
R8356 VSS.t20 VSS.n1932 25.542
R8357 VSS.t20 VSS.n1933 25.542
R8358 VSS.t20 VSS.n1934 25.542
R8359 VSS.t20 VSS.n1940 25.542
R8360 VSS.t20 VSS.n1941 25.542
R8361 VSS.t20 VSS.n1942 25.542
R8362 VSS.t20 VSS.n1943 25.542
R8363 VSS.t28 VSS.n1841 25.542
R8364 VSS.t28 VSS.n1842 25.542
R8365 VSS.t28 VSS.n1843 25.542
R8366 VSS.t28 VSS.n1844 25.542
R8367 VSS.t28 VSS.n1850 25.542
R8368 VSS.t28 VSS.n1851 25.542
R8369 VSS.t28 VSS.n1852 25.542
R8370 VSS.t28 VSS.n1853 25.542
R8371 VSS.t30 VSS.n1751 25.542
R8372 VSS.t30 VSS.n1752 25.542
R8373 VSS.t30 VSS.n1753 25.542
R8374 VSS.t30 VSS.n1754 25.542
R8375 VSS.t30 VSS.n1760 25.542
R8376 VSS.t30 VSS.n1761 25.542
R8377 VSS.t30 VSS.n1762 25.542
R8378 VSS.t30 VSS.n1763 25.542
R8379 VSS.t16 VSS.n1661 25.542
R8380 VSS.t16 VSS.n1662 25.542
R8381 VSS.t16 VSS.n1663 25.542
R8382 VSS.t16 VSS.n1664 25.542
R8383 VSS.t16 VSS.n1670 25.542
R8384 VSS.t16 VSS.n1671 25.542
R8385 VSS.t16 VSS.n1672 25.542
R8386 VSS.t16 VSS.n1673 25.542
R8387 VSS.t64 VSS.n6098 25.542
R8388 VSS.t64 VSS.n6096 25.542
R8389 VSS.t64 VSS.n6094 25.542
R8390 VSS.t64 VSS.n6092 25.542
R8391 VSS.t64 VSS.n6097 25.542
R8392 VSS.t64 VSS.n6095 25.542
R8393 VSS.t64 VSS.n6093 25.542
R8394 VSS.t64 VSS.n6091 25.542
R8395 VSS.t76 VSS.n5982 25.542
R8396 VSS.t76 VSS.n5980 25.542
R8397 VSS.t76 VSS.n5978 25.542
R8398 VSS.t76 VSS.n5976 25.542
R8399 VSS.t76 VSS.n5981 25.542
R8400 VSS.t76 VSS.n5979 25.542
R8401 VSS.t76 VSS.n5977 25.542
R8402 VSS.t76 VSS.n5975 25.542
R8403 VSS.t74 VSS.n5866 25.542
R8404 VSS.t74 VSS.n5864 25.542
R8405 VSS.t74 VSS.n5862 25.542
R8406 VSS.t74 VSS.n5860 25.542
R8407 VSS.t74 VSS.n5865 25.542
R8408 VSS.t74 VSS.n5863 25.542
R8409 VSS.t74 VSS.n5861 25.542
R8410 VSS.t74 VSS.n5859 25.542
R8411 VSS.n6992 VSS.t68 25.542
R8412 VSS.n6386 VSS.t68 25.542
R8413 VSS.n6985 VSS.t68 25.542
R8414 VSS.n6389 VSS.t68 25.542
R8415 VSS.n6943 VSS.t68 25.542
R8416 VSS.n6949 VSS.t68 25.542
R8417 VSS.n6396 VSS.t68 25.542
R8418 VSS.n6956 VSS.t68 25.542
R8419 VSS.t66 VSS.n6405 25.542
R8420 VSS.t66 VSS.n6406 25.542
R8421 VSS.t66 VSS.n6407 25.542
R8422 VSS.t66 VSS.n6408 25.542
R8423 VSS.t66 VSS.n6414 25.542
R8424 VSS.t66 VSS.n6415 25.542
R8425 VSS.t66 VSS.n6416 25.542
R8426 VSS.t66 VSS.n6417 25.542
R8427 VSS.t70 VSS.n6495 25.542
R8428 VSS.t70 VSS.n6496 25.542
R8429 VSS.t70 VSS.n6497 25.542
R8430 VSS.t70 VSS.n6498 25.542
R8431 VSS.t70 VSS.n6504 25.542
R8432 VSS.t70 VSS.n6505 25.542
R8433 VSS.t70 VSS.n6506 25.542
R8434 VSS.t70 VSS.n6507 25.542
R8435 VSS.t72 VSS.n6585 25.542
R8436 VSS.t72 VSS.n6586 25.542
R8437 VSS.t72 VSS.n6587 25.542
R8438 VSS.t72 VSS.n6588 25.542
R8439 VSS.t72 VSS.n6594 25.542
R8440 VSS.t72 VSS.n6595 25.542
R8441 VSS.t72 VSS.n6596 25.542
R8442 VSS.t72 VSS.n6597 25.542
R8443 VSS.t78 VSS.n17937 25.542
R8444 VSS.t78 VSS.n17926 25.542
R8445 VSS.t78 VSS.n17928 25.542
R8446 VSS.t78 VSS.n17930 25.542
R8447 VSS.t78 VSS.n17929 25.542
R8448 VSS.t78 VSS.n17931 25.542
R8449 VSS.n17643 VSS 23.829
R8450 VSS.n17980 VSS.n17977 23.644
R8451 VSS VSS.n18134 23.572
R8452 VSS.n18017 VSS.n17925 23.333
R8453 VSS.n392 VSS.n367 22.758
R8454 VSS.n420 VSS.n349 22.758
R8455 VSS.n18184 VSS.n18159 22.758
R8456 VSS.n18214 VSS.n18213 22.758
R8457 VSS.n17611 VSS 20.97
R8458 VSS.n18295 VSS 20
R8459 VSS.n408 VSS.n360 19.952
R8460 VSS.n408 VSS.n361 19.952
R8461 VSS.n18200 VSS.n18152 19.952
R8462 VSS.n18200 VSS.n18153 19.952
R8463 VSS.t78 VSS.n18016 19.67
R8464 VSS.n14655 VSS.n14651 19.504
R8465 VSS.n14669 VSS.n14665 19.504
R8466 VSS.n14683 VSS.n14679 19.504
R8467 VSS.n14697 VSS.n14693 19.504
R8468 VSS.n14711 VSS.n14707 19.504
R8469 VSS.n14729 VSS.n14721 19.504
R8470 VSS.n14747 VSS.n14743 19.504
R8471 VSS.n14761 VSS.n14757 19.504
R8472 VSS.n14775 VSS.n14771 19.504
R8473 VSS.n14789 VSS.n14785 19.504
R8474 VSS.n14807 VSS.n14799 19.504
R8475 VSS.n15155 VSS.n15151 19.504
R8476 VSS.n15169 VSS.n15165 19.504
R8477 VSS.n15183 VSS.n15179 19.504
R8478 VSS.n15197 VSS.n15193 19.504
R8479 VSS.n15211 VSS.n15207 19.504
R8480 VSS.n15229 VSS.n15221 19.504
R8481 VSS.n15247 VSS.n15243 19.504
R8482 VSS.n15261 VSS.n15257 19.504
R8483 VSS.n15275 VSS.n15271 19.504
R8484 VSS.n15289 VSS.n15285 19.504
R8485 VSS.n15307 VSS.n15299 19.504
R8486 VSS.n14911 VSS.n14907 19.504
R8487 VSS.n14925 VSS.n14921 19.504
R8488 VSS.n14939 VSS.n14935 19.504
R8489 VSS.n14953 VSS.n14949 19.504
R8490 VSS.n14967 VSS.n14963 19.504
R8491 VSS.n14985 VSS.n14977 19.504
R8492 VSS.n15003 VSS.n14999 19.504
R8493 VSS.n15017 VSS.n15013 19.504
R8494 VSS.n15031 VSS.n15027 19.504
R8495 VSS.n15045 VSS.n15041 19.504
R8496 VSS.n15063 VSS.n15055 19.504
R8497 VSS.n15643 VSS.n15639 19.504
R8498 VSS.n15657 VSS.n15653 19.504
R8499 VSS.n15671 VSS.n15667 19.504
R8500 VSS.n15685 VSS.n15681 19.504
R8501 VSS.n15699 VSS.n15695 19.504
R8502 VSS.n15717 VSS.n15709 19.504
R8503 VSS.n15735 VSS.n15731 19.504
R8504 VSS.n15749 VSS.n15745 19.504
R8505 VSS.n15763 VSS.n15759 19.504
R8506 VSS.n15777 VSS.n15773 19.504
R8507 VSS.n15795 VSS.n15787 19.504
R8508 VSS.n15399 VSS.n15395 19.504
R8509 VSS.n15413 VSS.n15409 19.504
R8510 VSS.n15427 VSS.n15423 19.504
R8511 VSS.n15441 VSS.n15437 19.504
R8512 VSS.n15455 VSS.n15451 19.504
R8513 VSS.n15473 VSS.n15465 19.504
R8514 VSS.n15491 VSS.n15487 19.504
R8515 VSS.n15505 VSS.n15501 19.504
R8516 VSS.n15519 VSS.n15515 19.504
R8517 VSS.n15533 VSS.n15529 19.504
R8518 VSS.n15551 VSS.n15543 19.504
R8519 VSS.n16131 VSS.n16127 19.504
R8520 VSS.n16145 VSS.n16141 19.504
R8521 VSS.n16159 VSS.n16155 19.504
R8522 VSS.n16173 VSS.n16169 19.504
R8523 VSS.n16187 VSS.n16183 19.504
R8524 VSS.n16205 VSS.n16197 19.504
R8525 VSS.n16223 VSS.n16219 19.504
R8526 VSS.n16237 VSS.n16233 19.504
R8527 VSS.n16251 VSS.n16247 19.504
R8528 VSS.n16265 VSS.n16261 19.504
R8529 VSS.n16283 VSS.n16275 19.504
R8530 VSS.n15887 VSS.n15883 19.504
R8531 VSS.n15901 VSS.n15897 19.504
R8532 VSS.n15915 VSS.n15911 19.504
R8533 VSS.n15929 VSS.n15925 19.504
R8534 VSS.n15943 VSS.n15939 19.504
R8535 VSS.n15961 VSS.n15953 19.504
R8536 VSS.n15979 VSS.n15975 19.504
R8537 VSS.n15993 VSS.n15989 19.504
R8538 VSS.n16007 VSS.n16003 19.504
R8539 VSS.n16021 VSS.n16017 19.504
R8540 VSS.n16039 VSS.n16031 19.504
R8541 VSS.n16387 VSS.n16383 19.504
R8542 VSS.n16401 VSS.n16397 19.504
R8543 VSS.n16415 VSS.n16411 19.504
R8544 VSS.n16429 VSS.n16425 19.504
R8545 VSS.n16443 VSS.n16439 19.504
R8546 VSS.n16461 VSS.n16453 19.504
R8547 VSS.n16479 VSS.n16475 19.504
R8548 VSS.n16493 VSS.n16489 19.504
R8549 VSS.n16507 VSS.n16503 19.504
R8550 VSS.n16521 VSS.n16517 19.504
R8551 VSS.n16582 VSS.n16576 19.504
R8552 VSS.n10704 VSS.n10700 19.504
R8553 VSS.n10718 VSS.n10714 19.504
R8554 VSS.n10732 VSS.n10728 19.504
R8555 VSS.n10746 VSS.n10742 19.504
R8556 VSS.n10760 VSS.n10756 19.504
R8557 VSS.n10778 VSS.n10770 19.504
R8558 VSS.n10796 VSS.n10792 19.504
R8559 VSS.n10810 VSS.n10806 19.504
R8560 VSS.n10824 VSS.n10820 19.504
R8561 VSS.n10838 VSS.n10834 19.504
R8562 VSS.n10856 VSS.n10848 19.504
R8563 VSS.n11204 VSS.n11200 19.504
R8564 VSS.n11218 VSS.n11214 19.504
R8565 VSS.n11232 VSS.n11228 19.504
R8566 VSS.n11246 VSS.n11242 19.504
R8567 VSS.n11260 VSS.n11256 19.504
R8568 VSS.n11278 VSS.n11270 19.504
R8569 VSS.n11296 VSS.n11292 19.504
R8570 VSS.n11310 VSS.n11306 19.504
R8571 VSS.n11324 VSS.n11320 19.504
R8572 VSS.n11338 VSS.n11334 19.504
R8573 VSS.n11356 VSS.n11348 19.504
R8574 VSS.n10960 VSS.n10956 19.504
R8575 VSS.n10974 VSS.n10970 19.504
R8576 VSS.n10988 VSS.n10984 19.504
R8577 VSS.n11002 VSS.n10998 19.504
R8578 VSS.n11016 VSS.n11012 19.504
R8579 VSS.n11034 VSS.n11026 19.504
R8580 VSS.n11052 VSS.n11048 19.504
R8581 VSS.n11066 VSS.n11062 19.504
R8582 VSS.n11080 VSS.n11076 19.504
R8583 VSS.n11094 VSS.n11090 19.504
R8584 VSS.n11112 VSS.n11104 19.504
R8585 VSS.n11692 VSS.n11688 19.504
R8586 VSS.n11706 VSS.n11702 19.504
R8587 VSS.n11720 VSS.n11716 19.504
R8588 VSS.n11734 VSS.n11730 19.504
R8589 VSS.n11748 VSS.n11744 19.504
R8590 VSS.n11766 VSS.n11758 19.504
R8591 VSS.n11784 VSS.n11780 19.504
R8592 VSS.n11798 VSS.n11794 19.504
R8593 VSS.n11812 VSS.n11808 19.504
R8594 VSS.n11826 VSS.n11822 19.504
R8595 VSS.n11844 VSS.n11836 19.504
R8596 VSS.n11448 VSS.n11444 19.504
R8597 VSS.n11462 VSS.n11458 19.504
R8598 VSS.n11476 VSS.n11472 19.504
R8599 VSS.n11490 VSS.n11486 19.504
R8600 VSS.n11504 VSS.n11500 19.504
R8601 VSS.n11522 VSS.n11514 19.504
R8602 VSS.n11540 VSS.n11536 19.504
R8603 VSS.n11554 VSS.n11550 19.504
R8604 VSS.n11568 VSS.n11564 19.504
R8605 VSS.n11582 VSS.n11578 19.504
R8606 VSS.n11600 VSS.n11592 19.504
R8607 VSS.n12180 VSS.n12176 19.504
R8608 VSS.n12194 VSS.n12190 19.504
R8609 VSS.n12208 VSS.n12204 19.504
R8610 VSS.n12222 VSS.n12218 19.504
R8611 VSS.n12236 VSS.n12232 19.504
R8612 VSS.n12254 VSS.n12246 19.504
R8613 VSS.n12272 VSS.n12268 19.504
R8614 VSS.n12286 VSS.n12282 19.504
R8615 VSS.n12300 VSS.n12296 19.504
R8616 VSS.n12314 VSS.n12310 19.504
R8617 VSS.n12332 VSS.n12324 19.504
R8618 VSS.n11936 VSS.n11932 19.504
R8619 VSS.n11950 VSS.n11946 19.504
R8620 VSS.n11964 VSS.n11960 19.504
R8621 VSS.n11978 VSS.n11974 19.504
R8622 VSS.n11992 VSS.n11988 19.504
R8623 VSS.n12010 VSS.n12002 19.504
R8624 VSS.n12028 VSS.n12024 19.504
R8625 VSS.n12042 VSS.n12038 19.504
R8626 VSS.n12056 VSS.n12052 19.504
R8627 VSS.n12070 VSS.n12066 19.504
R8628 VSS.n12088 VSS.n12080 19.504
R8629 VSS.n12436 VSS.n12432 19.504
R8630 VSS.n12450 VSS.n12446 19.504
R8631 VSS.n12464 VSS.n12460 19.504
R8632 VSS.n12478 VSS.n12474 19.504
R8633 VSS.n12492 VSS.n12488 19.504
R8634 VSS.n12510 VSS.n12502 19.504
R8635 VSS.n12528 VSS.n12524 19.504
R8636 VSS.n12542 VSS.n12538 19.504
R8637 VSS.n12556 VSS.n12552 19.504
R8638 VSS.n12570 VSS.n12566 19.504
R8639 VSS.n12631 VSS.n12625 19.504
R8640 VSS.n7272 VSS.n7268 19.504
R8641 VSS.n7286 VSS.n7282 19.504
R8642 VSS.n7300 VSS.n7296 19.504
R8643 VSS.n7314 VSS.n7310 19.504
R8644 VSS.n7328 VSS.n7324 19.504
R8645 VSS.n7346 VSS.n7338 19.504
R8646 VSS.n7364 VSS.n7360 19.504
R8647 VSS.n7378 VSS.n7374 19.504
R8648 VSS.n7392 VSS.n7388 19.504
R8649 VSS.n7406 VSS.n7402 19.504
R8650 VSS.n7424 VSS.n7416 19.504
R8651 VSS.n7772 VSS.n7768 19.504
R8652 VSS.n7786 VSS.n7782 19.504
R8653 VSS.n7800 VSS.n7796 19.504
R8654 VSS.n7814 VSS.n7810 19.504
R8655 VSS.n7828 VSS.n7824 19.504
R8656 VSS.n7846 VSS.n7838 19.504
R8657 VSS.n7864 VSS.n7860 19.504
R8658 VSS.n7878 VSS.n7874 19.504
R8659 VSS.n7892 VSS.n7888 19.504
R8660 VSS.n7906 VSS.n7902 19.504
R8661 VSS.n7924 VSS.n7916 19.504
R8662 VSS.n7528 VSS.n7524 19.504
R8663 VSS.n7542 VSS.n7538 19.504
R8664 VSS.n7556 VSS.n7552 19.504
R8665 VSS.n7570 VSS.n7566 19.504
R8666 VSS.n7584 VSS.n7580 19.504
R8667 VSS.n7602 VSS.n7594 19.504
R8668 VSS.n7620 VSS.n7616 19.504
R8669 VSS.n7634 VSS.n7630 19.504
R8670 VSS.n7648 VSS.n7644 19.504
R8671 VSS.n7662 VSS.n7658 19.504
R8672 VSS.n7680 VSS.n7672 19.504
R8673 VSS.n8260 VSS.n8256 19.504
R8674 VSS.n8274 VSS.n8270 19.504
R8675 VSS.n8288 VSS.n8284 19.504
R8676 VSS.n8302 VSS.n8298 19.504
R8677 VSS.n8316 VSS.n8312 19.504
R8678 VSS.n8334 VSS.n8326 19.504
R8679 VSS.n8352 VSS.n8348 19.504
R8680 VSS.n8366 VSS.n8362 19.504
R8681 VSS.n8380 VSS.n8376 19.504
R8682 VSS.n8394 VSS.n8390 19.504
R8683 VSS.n8412 VSS.n8404 19.504
R8684 VSS.n8016 VSS.n8012 19.504
R8685 VSS.n8030 VSS.n8026 19.504
R8686 VSS.n8044 VSS.n8040 19.504
R8687 VSS.n8058 VSS.n8054 19.504
R8688 VSS.n8072 VSS.n8068 19.504
R8689 VSS.n8090 VSS.n8082 19.504
R8690 VSS.n8108 VSS.n8104 19.504
R8691 VSS.n8122 VSS.n8118 19.504
R8692 VSS.n8136 VSS.n8132 19.504
R8693 VSS.n8150 VSS.n8146 19.504
R8694 VSS.n8168 VSS.n8160 19.504
R8695 VSS.n8748 VSS.n8744 19.504
R8696 VSS.n8762 VSS.n8758 19.504
R8697 VSS.n8776 VSS.n8772 19.504
R8698 VSS.n8790 VSS.n8786 19.504
R8699 VSS.n8804 VSS.n8800 19.504
R8700 VSS.n8822 VSS.n8814 19.504
R8701 VSS.n8840 VSS.n8836 19.504
R8702 VSS.n8854 VSS.n8850 19.504
R8703 VSS.n8868 VSS.n8864 19.504
R8704 VSS.n8882 VSS.n8878 19.504
R8705 VSS.n8900 VSS.n8892 19.504
R8706 VSS.n8504 VSS.n8500 19.504
R8707 VSS.n8518 VSS.n8514 19.504
R8708 VSS.n8532 VSS.n8528 19.504
R8709 VSS.n8546 VSS.n8542 19.504
R8710 VSS.n8560 VSS.n8556 19.504
R8711 VSS.n8578 VSS.n8570 19.504
R8712 VSS.n8596 VSS.n8592 19.504
R8713 VSS.n8610 VSS.n8606 19.504
R8714 VSS.n8624 VSS.n8620 19.504
R8715 VSS.n8638 VSS.n8634 19.504
R8716 VSS.n8656 VSS.n8648 19.504
R8717 VSS.n9004 VSS.n9000 19.504
R8718 VSS.n9018 VSS.n9014 19.504
R8719 VSS.n9032 VSS.n9028 19.504
R8720 VSS.n9046 VSS.n9042 19.504
R8721 VSS.n9060 VSS.n9056 19.504
R8722 VSS.n9078 VSS.n9070 19.504
R8723 VSS.n9096 VSS.n9092 19.504
R8724 VSS.n9110 VSS.n9106 19.504
R8725 VSS.n9124 VSS.n9120 19.504
R8726 VSS.n9138 VSS.n9134 19.504
R8727 VSS.n9199 VSS.n9193 19.504
R8728 VSS.n5140 VSS.n1584 19.504
R8729 VSS.n5148 VSS.n1577 19.504
R8730 VSS.n5159 VSS.n1571 19.504
R8731 VSS.n5163 VSS.n1565 19.504
R8732 VSS.n5175 VSS.n1563 19.504
R8733 VSS.n5183 VSS.n1556 19.504
R8734 VSS.n5194 VSS.n1550 19.504
R8735 VSS.n5198 VSS.n1544 19.504
R8736 VSS.n5210 VSS.n1542 19.504
R8737 VSS.n5218 VSS.n1534 19.504
R8738 VSS.n1535 VSS.n1529 19.504
R8739 VSS.n5403 VSS.n1526 19.504
R8740 VSS.n5499 VSS.n1443 19.504
R8741 VSS.n5507 VSS.n1436 19.504
R8742 VSS.n5518 VSS.n1430 19.504
R8743 VSS.n5522 VSS.n1424 19.504
R8744 VSS.n5534 VSS.n1422 19.504
R8745 VSS.n5542 VSS.n1415 19.504
R8746 VSS.n5553 VSS.n1409 19.504
R8747 VSS.n5557 VSS.n1403 19.504
R8748 VSS.n5569 VSS.n1401 19.504
R8749 VSS.n5577 VSS.n1393 19.504
R8750 VSS.n1394 VSS.n1388 19.504
R8751 VSS.n5611 VSS.n1385 19.504
R8752 VSS.n5398 VSS.n5236 19.504
R8753 VSS.n5386 VSS.n5240 19.504
R8754 VSS.n5379 VSS.n5249 19.504
R8755 VSS.n5375 VSS.n5253 19.504
R8756 VSS.n5363 VSS.n5260 19.504
R8757 VSS.n5356 VSS.n5268 19.504
R8758 VSS.n5352 VSS.n5272 19.504
R8759 VSS.n5340 VSS.n5279 19.504
R8760 VSS.n5333 VSS.n5287 19.504
R8761 VSS.n5329 VSS.n5291 19.504
R8762 VSS.n5317 VSS.n5298 19.504
R8763 VSS.n5310 VSS.n5307 19.504
R8764 VSS.n785 VSS.n780 19.504
R8765 VSS.n793 VSS.n773 19.504
R8766 VSS.n804 VSS.n767 19.504
R8767 VSS.n808 VSS.n761 19.504
R8768 VSS.n820 VSS.n759 19.504
R8769 VSS.n828 VSS.n752 19.504
R8770 VSS.n839 VSS.n746 19.504
R8771 VSS.n843 VSS.n740 19.504
R8772 VSS.n855 VSS.n738 19.504
R8773 VSS.n863 VSS.n731 19.504
R8774 VSS.n874 VSS.n724 19.504
R8775 VSS.n879 VSS.n878 19.504
R8776 VSS.n5606 VSS.n5595 19.504
R8777 VSS.n5781 VSS.n523 19.504
R8778 VSS.n5777 VSS.n527 19.504
R8779 VSS.n5765 VSS.n534 19.504
R8780 VSS.n5758 VSS.n542 19.504
R8781 VSS.n5754 VSS.n546 19.504
R8782 VSS.n5742 VSS.n553 19.504
R8783 VSS.n5735 VSS.n561 19.504
R8784 VSS.n5731 VSS.n565 19.504
R8785 VSS.n5719 VSS.n572 19.504
R8786 VSS.n5712 VSS.n580 19.504
R8787 VSS.n5708 VSS.n584 19.504
R8788 VSS.n920 VSS.n710 19.504
R8789 VSS.n932 VSS.n708 19.504
R8790 VSS.n940 VSS.n701 19.504
R8791 VSS.n951 VSS.n695 19.504
R8792 VSS.n955 VSS.n689 19.504
R8793 VSS.n967 VSS.n687 19.504
R8794 VSS.n975 VSS.n680 19.504
R8795 VSS.n986 VSS.n674 19.504
R8796 VSS.n990 VSS.n668 19.504
R8797 VSS.n1002 VSS.n666 19.504
R8798 VSS.n1010 VSS.n659 19.504
R8799 VSS.n1267 VSS.n654 19.504
R8800 VSS.n1258 VSS.n1023 19.504
R8801 VSS.n1254 VSS.n1027 19.504
R8802 VSS.n1242 VSS.n1034 19.504
R8803 VSS.n1235 VSS.n1042 19.504
R8804 VSS.n1231 VSS.n1046 19.504
R8805 VSS.n1219 VSS.n1053 19.504
R8806 VSS.n1212 VSS.n1061 19.504
R8807 VSS.n1208 VSS.n1065 19.504
R8808 VSS.n1196 VSS.n1072 19.504
R8809 VSS.n1189 VSS.n1080 19.504
R8810 VSS.n1185 VSS.n1084 19.504
R8811 VSS.n1173 VSS.n1091 19.504
R8812 VSS.n3805 VSS.n3450 19.504
R8813 VSS.n3801 VSS.n3456 19.504
R8814 VSS.n3789 VSS.n3464 19.504
R8815 VSS.n3782 VSS.n3472 19.504
R8816 VSS.n3778 VSS.n3476 19.504
R8817 VSS.n3766 VSS.n3483 19.504
R8818 VSS.n3759 VSS.n3491 19.504
R8819 VSS.n3755 VSS.n3495 19.504
R8820 VSS.n3743 VSS.n3502 19.504
R8821 VSS.n3736 VSS.n3510 19.504
R8822 VSS.n3732 VSS.n3514 19.504
R8823 VSS.n3720 VSS.n3521 19.504
R8824 VSS.n3962 VSS.n3380 19.504
R8825 VSS.n3974 VSS.n3378 19.504
R8826 VSS.n3982 VSS.n3371 19.504
R8827 VSS.n3993 VSS.n3365 19.504
R8828 VSS.n3997 VSS.n3359 19.504
R8829 VSS.n4009 VSS.n3357 19.504
R8830 VSS.n4017 VSS.n3350 19.504
R8831 VSS.n4028 VSS.n3344 19.504
R8832 VSS.n4032 VSS.n3338 19.504
R8833 VSS.n4044 VSS.n3336 19.504
R8834 VSS.n4052 VSS.n3329 19.504
R8835 VSS.n4418 VSS.n3324 19.504
R8836 VSS.n3712 VSS.n3562 19.504
R8837 VSS.n3708 VSS.n3569 19.504
R8838 VSS.n3696 VSS.n3576 19.504
R8839 VSS.n3689 VSS.n3584 19.504
R8840 VSS.n3685 VSS.n3588 19.504
R8841 VSS.n3673 VSS.n3595 19.504
R8842 VSS.n3666 VSS.n3603 19.504
R8843 VSS.n3662 VSS.n3607 19.504
R8844 VSS.n3650 VSS.n3614 19.504
R8845 VSS.n3643 VSS.n3622 19.504
R8846 VSS.n3639 VSS.n3626 19.504
R8847 VSS.n3957 VSS.n3387 19.504
R8848 VSS.n4316 VSS.n4174 19.504
R8849 VSS.n4312 VSS.n4181 19.504
R8850 VSS.n4300 VSS.n4188 19.504
R8851 VSS.n4293 VSS.n4196 19.504
R8852 VSS.n4289 VSS.n4200 19.504
R8853 VSS.n4277 VSS.n4207 19.504
R8854 VSS.n4270 VSS.n4215 19.504
R8855 VSS.n4266 VSS.n4219 19.504
R8856 VSS.n4254 VSS.n4226 19.504
R8857 VSS.n4247 VSS.n4234 19.504
R8858 VSS.n4243 VSS.n3225 19.504
R8859 VSS.n4531 VSS.n3226 19.504
R8860 VSS.n4409 VSS.n4065 19.504
R8861 VSS.n4405 VSS.n4069 19.504
R8862 VSS.n4393 VSS.n4076 19.504
R8863 VSS.n4386 VSS.n4084 19.504
R8864 VSS.n4382 VSS.n4088 19.504
R8865 VSS.n4370 VSS.n4095 19.504
R8866 VSS.n4363 VSS.n4103 19.504
R8867 VSS.n4359 VSS.n4107 19.504
R8868 VSS.n4347 VSS.n4114 19.504
R8869 VSS.n4340 VSS.n4122 19.504
R8870 VSS.n4336 VSS.n4126 19.504
R8871 VSS.n4324 VSS.n4133 19.504
R8872 VSS.n5018 VSS.n4653 19.504
R8873 VSS.n5014 VSS.n4659 19.504
R8874 VSS.n5002 VSS.n4666 19.504
R8875 VSS.n4995 VSS.n4674 19.504
R8876 VSS.n4991 VSS.n4678 19.504
R8877 VSS.n4979 VSS.n4685 19.504
R8878 VSS.n4972 VSS.n4693 19.504
R8879 VSS.n4968 VSS.n4697 19.504
R8880 VSS.n4956 VSS.n4704 19.504
R8881 VSS.n4949 VSS.n4712 19.504
R8882 VSS.n4945 VSS.n4716 19.504
R8883 VSS.n4933 VSS.n4723 19.504
R8884 VSS.n4548 VSS.n3215 19.504
R8885 VSS.n4559 VSS.n3209 19.504
R8886 VSS.n4563 VSS.n3203 19.504
R8887 VSS.n4575 VSS.n3201 19.504
R8888 VSS.n4583 VSS.n3194 19.504
R8889 VSS.n4594 VSS.n3188 19.504
R8890 VSS.n4598 VSS.n3182 19.504
R8891 VSS.n4610 VSS.n3180 19.504
R8892 VSS.n4618 VSS.n3173 19.504
R8893 VSS.n4629 VSS.n3167 19.504
R8894 VSS.n4633 VSS.n3161 19.504
R8895 VSS.n4645 VSS.n3159 19.504
R8896 VSS.n4925 VSS.n4764 19.504
R8897 VSS.n4921 VSS.n4771 19.504
R8898 VSS.n4909 VSS.n4778 19.504
R8899 VSS.n4902 VSS.n4786 19.504
R8900 VSS.n4898 VSS.n4790 19.504
R8901 VSS.n4886 VSS.n4797 19.504
R8902 VSS.n4879 VSS.n4805 19.504
R8903 VSS.n4875 VSS.n4809 19.504
R8904 VSS.n4863 VSS.n4816 19.504
R8905 VSS.n4856 VSS.n4824 19.504
R8906 VSS.n4852 VSS.n4828 19.504
R8907 VSS.n4840 VSS.n4835 19.504
R8908 VSS.t6 VSS.n17550 19.3
R8909 VSS.t2 VSS.n17382 19.3
R8910 VSS.t4 VSS.n17214 19.3
R8911 VSS.t12 VSS.n17046 19.3
R8912 VSS.t14 VSS.n16878 19.3
R8913 VSS.t0 VSS.n16710 19.3
R8914 VSS.t56 VSS.n10515 19.3
R8915 VSS.t64 VSS.n6089 19.3
R8916 VSS.t76 VSS.n5973 19.3
R8917 VSS.t74 VSS.n5857 19.3
R8918 VSS.n6978 VSS.t68 19.3
R8919 VSS.t78 VSS.n17936 19.3
R8920 VSS.n385 VSS.n371 18.62
R8921 VSS.n428 VSS.n427 18.62
R8922 VSS.n18177 VSS.n18163 18.62
R8923 VSS.n18223 VSS.n18222 18.62
R8924 VSS.n14802 VSS.n14801 18.614
R8925 VSS.n15058 VSS.n15057 18.614
R8926 VSS.n15302 VSS.n15301 18.614
R8927 VSS.n15546 VSS.n15545 18.614
R8928 VSS.n15790 VSS.n15789 18.614
R8929 VSS.n16034 VSS.n16033 18.614
R8930 VSS.n16278 VSS.n16277 18.614
R8931 VSS.n10851 VSS.n10850 18.614
R8932 VSS.n11107 VSS.n11106 18.614
R8933 VSS.n11351 VSS.n11350 18.614
R8934 VSS.n11595 VSS.n11594 18.614
R8935 VSS.n11839 VSS.n11838 18.614
R8936 VSS.n12083 VSS.n12082 18.614
R8937 VSS.n12327 VSS.n12326 18.614
R8938 VSS.n7419 VSS.n7418 18.614
R8939 VSS.n7675 VSS.n7674 18.614
R8940 VSS.n7919 VSS.n7918 18.614
R8941 VSS.n8163 VSS.n8162 18.614
R8942 VSS.n8407 VSS.n8406 18.614
R8943 VSS.n8651 VSS.n8650 18.614
R8944 VSS.n8895 VSS.n8894 18.614
R8945 VSS.n1527 VSS.n1520 18.614
R8946 VSS.n5491 VSS.n1445 18.614
R8947 VSS.n1386 VSS.n1379 18.614
R8948 VSS.n5699 VSS.n592 18.614
R8949 VSS.n915 VSS.n717 18.614
R8950 VSS.n1271 VSS.n651 18.614
R8951 VSS.n3556 VSS.n3523 18.614
R8952 VSS.n3949 VSS.n3388 18.614
R8953 VSS.n4422 VSS.n3321 18.614
R8954 VSS.n4168 VSS.n4135 18.614
R8955 VSS.n4530 VSS.n4529 18.614
R8956 VSS.n5024 VSS.n3154 18.614
R8957 VSS.n4758 VSS.n4725 18.614
R8958 VSS.n378 VSS.n377 18.219
R8959 VSS.n436 VSS.n435 18.219
R8960 VSS.n18170 VSS.n18169 18.219
R8961 VSS.n18227 VSS.n18135 18.219
R8962 VSS.n14101 VSS 18.112
R8963 VSS.n14608 VSS.n14605 17.453
R8964 VSS.n10657 VSS.n10654 17.453
R8965 VSS.n7225 VSS.n7222 17.453
R8966 VSS.n1629 VSS.n1628 17.453
R8967 VSS.n3838 VSS.n3434 17.453
R8968 VSS.n17831 VSS.n17820 17.453
R8969 VSS.n17998 VSS.n17996 17.422
R8970 VSS.n16536 VSS.n16533 17.065
R8971 VSS.n12585 VSS.n12582 17.065
R8972 VSS.n9153 VSS.n9150 17.065
R8973 VSS.n1142 VSS.n1141 17.065
R8974 VSS.n5105 VSS.n5104 17.065
R8975 VSS.n17905 VSS.n17904 17.065
R8976 VSS.n14319 VSS.n14317 16.666
R8977 VSS.n14331 VSS.n14329 16.666
R8978 VSS.n14343 VSS.n14341 16.666
R8979 VSS.n14355 VSS.n14353 16.666
R8980 VSS.n14367 VSS.n14365 16.666
R8981 VSS.n14379 VSS.n14377 16.666
R8982 VSS.n14391 VSS.n14389 16.666
R8983 VSS.n14403 VSS.n14401 16.666
R8984 VSS.n14139 VSS.n14137 16.666
R8985 VSS.n14151 VSS.n14149 16.666
R8986 VSS.n14163 VSS.n14161 16.666
R8987 VSS.n14175 VSS.n14173 16.666
R8988 VSS.n14187 VSS.n14185 16.666
R8989 VSS.n14199 VSS.n14197 16.666
R8990 VSS.n14211 VSS.n14209 16.666
R8991 VSS.n14223 VSS.n14221 16.666
R8992 VSS.n17580 VSS.n17532 16.666
R8993 VSS.n17521 VSS.n17519 16.666
R8994 VSS.n17509 VSS.n17507 16.666
R8995 VSS.n17497 VSS.n17495 16.666
R8996 VSS.n17485 VSS.n17483 16.666
R8997 VSS.n17476 VSS.n17474 16.666
R8998 VSS.n17461 VSS.n17459 16.666
R8999 VSS.n17449 VSS.n17447 16.666
R9000 VSS.n17412 VSS.n17364 16.666
R9001 VSS.n17353 VSS.n17351 16.666
R9002 VSS.n17341 VSS.n17339 16.666
R9003 VSS.n17329 VSS.n17327 16.666
R9004 VSS.n17317 VSS.n17315 16.666
R9005 VSS.n17308 VSS.n17306 16.666
R9006 VSS.n17293 VSS.n17291 16.666
R9007 VSS.n17281 VSS.n17279 16.666
R9008 VSS.n17244 VSS.n17196 16.666
R9009 VSS.n17185 VSS.n17183 16.666
R9010 VSS.n17173 VSS.n17171 16.666
R9011 VSS.n17161 VSS.n17159 16.666
R9012 VSS.n17149 VSS.n17147 16.666
R9013 VSS.n17140 VSS.n17138 16.666
R9014 VSS.n17125 VSS.n17123 16.666
R9015 VSS.n17113 VSS.n17111 16.666
R9016 VSS.n17076 VSS.n17028 16.666
R9017 VSS.n17017 VSS.n17015 16.666
R9018 VSS.n17005 VSS.n17003 16.666
R9019 VSS.n16993 VSS.n16991 16.666
R9020 VSS.n16981 VSS.n16979 16.666
R9021 VSS.n16972 VSS.n16970 16.666
R9022 VSS.n16957 VSS.n16955 16.666
R9023 VSS.n16945 VSS.n16943 16.666
R9024 VSS.n16908 VSS.n16860 16.666
R9025 VSS.n16849 VSS.n16847 16.666
R9026 VSS.n16837 VSS.n16835 16.666
R9027 VSS.n16825 VSS.n16823 16.666
R9028 VSS.n16813 VSS.n16811 16.666
R9029 VSS.n16804 VSS.n16802 16.666
R9030 VSS.n16789 VSS.n16787 16.666
R9031 VSS.n16777 VSS.n16775 16.666
R9032 VSS.n16740 VSS.n16692 16.666
R9033 VSS.n16681 VSS.n16679 16.666
R9034 VSS.n16669 VSS.n16667 16.666
R9035 VSS.n16657 VSS.n16655 16.666
R9036 VSS.n16645 VSS.n16643 16.666
R9037 VSS.n16636 VSS.n16634 16.666
R9038 VSS.n16621 VSS.n16619 16.666
R9039 VSS.n16609 VSS.n16607 16.666
R9040 VSS.n13916 VSS.n13914 16.666
R9041 VSS.n13928 VSS.n13926 16.666
R9042 VSS.n13940 VSS.n13938 16.666
R9043 VSS.n13952 VSS.n13950 16.666
R9044 VSS.n13964 VSS.n13962 16.666
R9045 VSS.n13976 VSS.n13974 16.666
R9046 VSS.n13988 VSS.n13986 16.666
R9047 VSS.n14000 VSS.n13998 16.666
R9048 VSS.n13736 VSS.n13734 16.666
R9049 VSS.n13748 VSS.n13746 16.666
R9050 VSS.n13760 VSS.n13758 16.666
R9051 VSS.n13772 VSS.n13770 16.666
R9052 VSS.n13784 VSS.n13782 16.666
R9053 VSS.n13796 VSS.n13794 16.666
R9054 VSS.n13808 VSS.n13806 16.666
R9055 VSS.n13820 VSS.n13818 16.666
R9056 VSS.n13556 VSS.n13554 16.666
R9057 VSS.n13568 VSS.n13566 16.666
R9058 VSS.n13580 VSS.n13578 16.666
R9059 VSS.n13592 VSS.n13590 16.666
R9060 VSS.n13604 VSS.n13602 16.666
R9061 VSS.n13616 VSS.n13614 16.666
R9062 VSS.n13628 VSS.n13626 16.666
R9063 VSS.n13640 VSS.n13638 16.666
R9064 VSS.n13376 VSS.n13374 16.666
R9065 VSS.n13388 VSS.n13386 16.666
R9066 VSS.n13400 VSS.n13398 16.666
R9067 VSS.n13412 VSS.n13410 16.666
R9068 VSS.n13424 VSS.n13422 16.666
R9069 VSS.n13436 VSS.n13434 16.666
R9070 VSS.n13448 VSS.n13446 16.666
R9071 VSS.n13460 VSS.n13458 16.666
R9072 VSS.n13196 VSS.n13194 16.666
R9073 VSS.n13208 VSS.n13206 16.666
R9074 VSS.n13220 VSS.n13218 16.666
R9075 VSS.n13232 VSS.n13230 16.666
R9076 VSS.n13244 VSS.n13242 16.666
R9077 VSS.n13256 VSS.n13254 16.666
R9078 VSS.n13268 VSS.n13266 16.666
R9079 VSS.n13280 VSS.n13278 16.666
R9080 VSS.n13016 VSS.n13014 16.666
R9081 VSS.n13028 VSS.n13026 16.666
R9082 VSS.n13040 VSS.n13038 16.666
R9083 VSS.n13052 VSS.n13050 16.666
R9084 VSS.n13064 VSS.n13062 16.666
R9085 VSS.n13076 VSS.n13074 16.666
R9086 VSS.n13088 VSS.n13086 16.666
R9087 VSS.n13100 VSS.n13098 16.666
R9088 VSS.n12836 VSS.n12834 16.666
R9089 VSS.n12848 VSS.n12846 16.666
R9090 VSS.n12860 VSS.n12858 16.666
R9091 VSS.n12872 VSS.n12870 16.666
R9092 VSS.n12884 VSS.n12882 16.666
R9093 VSS.n12896 VSS.n12894 16.666
R9094 VSS.n12908 VSS.n12906 16.666
R9095 VSS.n12920 VSS.n12918 16.666
R9096 VSS.n12656 VSS.n12654 16.666
R9097 VSS.n12668 VSS.n12666 16.666
R9098 VSS.n12680 VSS.n12678 16.666
R9099 VSS.n12692 VSS.n12690 16.666
R9100 VSS.n12704 VSS.n12702 16.666
R9101 VSS.n12716 VSS.n12714 16.666
R9102 VSS.n12728 VSS.n12726 16.666
R9103 VSS.n12740 VSS.n12738 16.666
R9104 VSS.n9368 VSS.n9321 16.666
R9105 VSS.n9311 VSS.n9309 16.666
R9106 VSS.n9299 VSS.n9297 16.666
R9107 VSS.n9287 VSS.n9285 16.666
R9108 VSS.n9275 VSS.n9273 16.666
R9109 VSS.n9266 VSS.n9264 16.666
R9110 VSS.n9251 VSS.n9249 16.666
R9111 VSS.n9239 VSS.n9237 16.666
R9112 VSS.n9536 VSS.n9489 16.666
R9113 VSS.n9479 VSS.n9477 16.666
R9114 VSS.n9467 VSS.n9465 16.666
R9115 VSS.n9455 VSS.n9453 16.666
R9116 VSS.n9443 VSS.n9441 16.666
R9117 VSS.n9434 VSS.n9432 16.666
R9118 VSS.n9419 VSS.n9417 16.666
R9119 VSS.n9407 VSS.n9405 16.666
R9120 VSS.n9704 VSS.n9657 16.666
R9121 VSS.n9647 VSS.n9645 16.666
R9122 VSS.n9635 VSS.n9633 16.666
R9123 VSS.n9623 VSS.n9621 16.666
R9124 VSS.n9611 VSS.n9609 16.666
R9125 VSS.n9602 VSS.n9600 16.666
R9126 VSS.n9587 VSS.n9585 16.666
R9127 VSS.n9575 VSS.n9573 16.666
R9128 VSS.n9872 VSS.n9825 16.666
R9129 VSS.n9815 VSS.n9813 16.666
R9130 VSS.n9803 VSS.n9801 16.666
R9131 VSS.n9791 VSS.n9789 16.666
R9132 VSS.n9779 VSS.n9777 16.666
R9133 VSS.n9770 VSS.n9768 16.666
R9134 VSS.n9755 VSS.n9753 16.666
R9135 VSS.n9743 VSS.n9741 16.666
R9136 VSS.n10040 VSS.n9993 16.666
R9137 VSS.n9983 VSS.n9981 16.666
R9138 VSS.n9971 VSS.n9969 16.666
R9139 VSS.n9959 VSS.n9957 16.666
R9140 VSS.n9947 VSS.n9945 16.666
R9141 VSS.n9938 VSS.n9936 16.666
R9142 VSS.n9923 VSS.n9921 16.666
R9143 VSS.n9911 VSS.n9909 16.666
R9144 VSS.n10208 VSS.n10161 16.666
R9145 VSS.n10151 VSS.n10149 16.666
R9146 VSS.n10139 VSS.n10137 16.666
R9147 VSS.n10127 VSS.n10125 16.666
R9148 VSS.n10115 VSS.n10113 16.666
R9149 VSS.n10106 VSS.n10104 16.666
R9150 VSS.n10091 VSS.n10089 16.666
R9151 VSS.n10079 VSS.n10077 16.666
R9152 VSS.n10376 VSS.n10329 16.666
R9153 VSS.n10319 VSS.n10317 16.666
R9154 VSS.n10307 VSS.n10305 16.666
R9155 VSS.n10295 VSS.n10293 16.666
R9156 VSS.n10283 VSS.n10281 16.666
R9157 VSS.n10274 VSS.n10272 16.666
R9158 VSS.n10259 VSS.n10257 16.666
R9159 VSS.n10247 VSS.n10245 16.666
R9160 VSS.n10544 VSS.n10497 16.666
R9161 VSS.n10486 VSS.n10484 16.666
R9162 VSS.n10474 VSS.n10472 16.666
R9163 VSS.n10462 VSS.n10460 16.666
R9164 VSS.n10450 VSS.n10448 16.666
R9165 VSS.n10441 VSS.n10439 16.666
R9166 VSS.n10426 VSS.n10424 16.666
R9167 VSS.n10414 VSS.n10412 16.666
R9168 VSS.n2323 VSS.n2309 16.666
R9169 VSS.n2452 VSS.n2306 16.666
R9170 VSS.n2443 VSS.n2310 16.666
R9171 VSS.n2437 VSS.n2305 16.666
R9172 VSS.n2431 VSS.n2311 16.666
R9173 VSS.n2425 VSS.n2304 16.666
R9174 VSS.n2459 VSS.n2313 16.666
R9175 VSS.n2414 VSS.n2308 16.666
R9176 VSS.n2406 VSS.n2288 16.666
R9177 VSS.n2233 VSS.n2219 16.666
R9178 VSS.n2542 VSS.n2216 16.666
R9179 VSS.n2533 VSS.n2220 16.666
R9180 VSS.n2527 VSS.n2215 16.666
R9181 VSS.n2521 VSS.n2221 16.666
R9182 VSS.n2515 VSS.n2214 16.666
R9183 VSS.n2549 VSS.n2223 16.666
R9184 VSS.n2504 VSS.n2218 16.666
R9185 VSS.n2496 VSS.n2198 16.666
R9186 VSS.n2143 VSS.n2129 16.666
R9187 VSS.n2632 VSS.n2126 16.666
R9188 VSS.n2623 VSS.n2130 16.666
R9189 VSS.n2617 VSS.n2125 16.666
R9190 VSS.n2611 VSS.n2131 16.666
R9191 VSS.n2605 VSS.n2124 16.666
R9192 VSS.n2639 VSS.n2133 16.666
R9193 VSS.n2594 VSS.n2128 16.666
R9194 VSS.n2586 VSS.n2108 16.666
R9195 VSS.n2053 VSS.n2039 16.666
R9196 VSS.n2722 VSS.n2036 16.666
R9197 VSS.n2713 VSS.n2040 16.666
R9198 VSS.n2707 VSS.n2035 16.666
R9199 VSS.n2701 VSS.n2041 16.666
R9200 VSS.n2695 VSS.n2034 16.666
R9201 VSS.n2729 VSS.n2043 16.666
R9202 VSS.n2684 VSS.n2038 16.666
R9203 VSS.n2676 VSS.n2018 16.666
R9204 VSS.n1963 VSS.n1949 16.666
R9205 VSS.n2812 VSS.n1946 16.666
R9206 VSS.n2803 VSS.n1950 16.666
R9207 VSS.n2797 VSS.n1945 16.666
R9208 VSS.n2791 VSS.n1951 16.666
R9209 VSS.n2785 VSS.n1944 16.666
R9210 VSS.n2819 VSS.n1953 16.666
R9211 VSS.n2774 VSS.n1948 16.666
R9212 VSS.n2766 VSS.n1928 16.666
R9213 VSS.n1873 VSS.n1859 16.666
R9214 VSS.n2902 VSS.n1856 16.666
R9215 VSS.n2893 VSS.n1860 16.666
R9216 VSS.n2887 VSS.n1855 16.666
R9217 VSS.n2881 VSS.n1861 16.666
R9218 VSS.n2875 VSS.n1854 16.666
R9219 VSS.n2909 VSS.n1863 16.666
R9220 VSS.n2864 VSS.n1858 16.666
R9221 VSS.n2856 VSS.n1838 16.666
R9222 VSS.n1783 VSS.n1769 16.666
R9223 VSS.n2992 VSS.n1766 16.666
R9224 VSS.n2983 VSS.n1770 16.666
R9225 VSS.n2977 VSS.n1765 16.666
R9226 VSS.n2971 VSS.n1771 16.666
R9227 VSS.n2965 VSS.n1764 16.666
R9228 VSS.n2999 VSS.n1773 16.666
R9229 VSS.n2954 VSS.n1768 16.666
R9230 VSS.n2946 VSS.n1748 16.666
R9231 VSS.n1693 VSS.n1679 16.666
R9232 VSS.n3082 VSS.n1676 16.666
R9233 VSS.n3073 VSS.n1680 16.666
R9234 VSS.n3067 VSS.n1675 16.666
R9235 VSS.n3061 VSS.n1681 16.666
R9236 VSS.n3055 VSS.n1674 16.666
R9237 VSS.n3089 VSS.n1683 16.666
R9238 VSS.n3044 VSS.n1678 16.666
R9239 VSS.n3036 VSS.n1658 16.666
R9240 VSS.n6126 VSS.n6077 16.666
R9241 VSS.n6134 VSS.n6081 16.666
R9242 VSS.n6142 VSS.n6080 16.666
R9243 VSS.n6150 VSS.n6082 16.666
R9244 VSS.n6158 VSS.n6079 16.666
R9245 VSS.n6166 VSS.n6083 16.666
R9246 VSS.n6174 VSS.n6078 16.666
R9247 VSS.n6182 VSS.n6084 16.666
R9248 VSS.n6010 VSS.n5961 16.666
R9249 VSS.n6018 VSS.n5965 16.666
R9250 VSS.n6026 VSS.n5964 16.666
R9251 VSS.n6034 VSS.n5966 16.666
R9252 VSS.n6042 VSS.n5963 16.666
R9253 VSS.n6050 VSS.n5967 16.666
R9254 VSS.n6058 VSS.n5962 16.666
R9255 VSS.n6066 VSS.n5968 16.666
R9256 VSS.n5894 VSS.n5845 16.666
R9257 VSS.n5902 VSS.n5849 16.666
R9258 VSS.n5910 VSS.n5848 16.666
R9259 VSS.n5918 VSS.n5850 16.666
R9260 VSS.n5926 VSS.n5847 16.666
R9261 VSS.n5934 VSS.n5851 16.666
R9262 VSS.n5942 VSS.n5846 16.666
R9263 VSS.n5950 VSS.n5852 16.666
R9264 VSS.n7042 VSS.n5789 16.666
R9265 VSS.n7036 VSS.n5790 16.666
R9266 VSS.n7030 VSS.n5795 16.666
R9267 VSS.n7024 VSS.n5801 16.666
R9268 VSS.n7018 VSS.n5807 16.666
R9269 VSS.n7012 VSS.n5813 16.666
R9270 VSS.n7006 VSS.n5818 16.666
R9271 VSS.n7000 VSS.n5825 16.666
R9272 VSS.n6851 VSS.n6437 16.666
R9273 VSS.n6925 VSS.n6423 16.666
R9274 VSS.n6916 VSS.n6420 16.666
R9275 VSS.n6910 VSS.n6424 16.666
R9276 VSS.n6904 VSS.n6419 16.666
R9277 VSS.n6898 VSS.n6425 16.666
R9278 VSS.n6892 VSS.n6418 16.666
R9279 VSS.n6933 VSS.n6427 16.666
R9280 VSS.n6761 VSS.n6527 16.666
R9281 VSS.n6835 VSS.n6513 16.666
R9282 VSS.n6826 VSS.n6510 16.666
R9283 VSS.n6820 VSS.n6514 16.666
R9284 VSS.n6814 VSS.n6509 16.666
R9285 VSS.n6808 VSS.n6515 16.666
R9286 VSS.n6802 VSS.n6508 16.666
R9287 VSS.n6843 VSS.n6517 16.666
R9288 VSS.n6671 VSS.n6617 16.666
R9289 VSS.n6745 VSS.n6603 16.666
R9290 VSS.n6736 VSS.n6600 16.666
R9291 VSS.n6730 VSS.n6604 16.666
R9292 VSS.n6724 VSS.n6599 16.666
R9293 VSS.n6718 VSS.n6605 16.666
R9294 VSS.n6712 VSS.n6598 16.666
R9295 VSS.n6753 VSS.n6607 16.666
R9296 VSS.n379 VSS.n371 16.551
R9297 VSS.n427 VSS.n344 16.551
R9298 VSS.n18171 VSS.n18163 16.551
R9299 VSS.n18224 VSS.n18223 16.551
R9300 VSS.n14477 VSS.n14475 16
R9301 VSS.n14475 VSS.n14474 16
R9302 VSS.n14474 VSS.n14473 16
R9303 VSS.n14473 VSS.n14472 16
R9304 VSS.n14472 VSS.n14471 16
R9305 VSS.n14471 VSS.n14470 16
R9306 VSS.n14470 VSS.n14469 16
R9307 VSS.n14469 VSS.n14468 16
R9308 VSS.n14467 VSS.n14466 16
R9309 VSS.n14310 VSS.n14308 16
R9310 VSS.n14308 VSS.n14307 16
R9311 VSS.n14307 VSS.n14306 16
R9312 VSS.n14306 VSS.n14305 16
R9313 VSS.n14305 VSS.n14304 16
R9314 VSS.n14304 VSS.n14303 16
R9315 VSS.n14303 VSS.n14302 16
R9316 VSS.n14302 VSS.n14301 16
R9317 VSS.n14297 VSS.n14295 16
R9318 VSS.n14295 VSS.n14294 16
R9319 VSS.n14294 VSS.n14293 16
R9320 VSS.n14293 VSS.n14292 16
R9321 VSS.n14292 VSS.n14291 16
R9322 VSS.n14291 VSS.n14290 16
R9323 VSS.n14290 VSS.n14289 16
R9324 VSS.n14289 VSS.n14288 16
R9325 VSS.n14287 VSS.n14286 16
R9326 VSS.n14131 VSS.n14129 16
R9327 VSS.n14129 VSS.n14128 16
R9328 VSS.n14128 VSS.n14127 16
R9329 VSS.n14127 VSS.n14126 16
R9330 VSS.n14126 VSS.n14125 16
R9331 VSS.n14125 VSS.n14124 16
R9332 VSS.n14124 VSS.n14123 16
R9333 VSS.n14123 VSS.n14122 16
R9334 VSS.n14490 VSS.n14489 16
R9335 VSS.n14489 VSS.n14488 16
R9336 VSS.n14488 VSS.n14487 16
R9337 VSS.n14487 VSS.n14486 16
R9338 VSS.n14486 VSS.n14485 16
R9339 VSS.n14485 VSS.n14484 16
R9340 VSS.n14484 VSS.n14483 16
R9341 VSS.n14483 VSS.n14482 16
R9342 VSS.n14481 VSS.n14480 16
R9343 VSS.n17595 VSS.n17594 16
R9344 VSS.n17594 VSS.n17593 16
R9345 VSS.n17593 VSS.n17592 16
R9346 VSS.n17592 VSS.n17591 16
R9347 VSS.n17591 VSS.n17590 16
R9348 VSS.n17590 VSS.n17589 16
R9349 VSS.n17589 VSS.n17588 16
R9350 VSS.n17588 VSS.n17587 16
R9351 VSS.n14502 VSS.n14501 16
R9352 VSS.n14501 VSS.n14500 16
R9353 VSS.n14500 VSS.n14499 16
R9354 VSS.n14499 VSS.n14498 16
R9355 VSS.n14498 VSS.n14497 16
R9356 VSS.n14497 VSS.n14496 16
R9357 VSS.n14496 VSS.n14495 16
R9358 VSS.n14495 VSS.n14494 16
R9359 VSS.n14493 VSS.n14492 16
R9360 VSS.n17427 VSS.n17426 16
R9361 VSS.n17426 VSS.n17425 16
R9362 VSS.n17425 VSS.n17424 16
R9363 VSS.n17424 VSS.n17423 16
R9364 VSS.n17423 VSS.n17422 16
R9365 VSS.n17422 VSS.n17421 16
R9366 VSS.n17421 VSS.n17420 16
R9367 VSS.n17420 VSS.n17419 16
R9368 VSS.n14514 VSS.n14513 16
R9369 VSS.n14513 VSS.n14512 16
R9370 VSS.n14512 VSS.n14511 16
R9371 VSS.n14511 VSS.n14510 16
R9372 VSS.n14510 VSS.n14509 16
R9373 VSS.n14509 VSS.n14508 16
R9374 VSS.n14508 VSS.n14507 16
R9375 VSS.n14507 VSS.n14506 16
R9376 VSS.n14505 VSS.n14504 16
R9377 VSS.n17259 VSS.n17258 16
R9378 VSS.n17258 VSS.n17257 16
R9379 VSS.n17257 VSS.n17256 16
R9380 VSS.n17256 VSS.n17255 16
R9381 VSS.n17255 VSS.n17254 16
R9382 VSS.n17254 VSS.n17253 16
R9383 VSS.n17253 VSS.n17252 16
R9384 VSS.n17252 VSS.n17251 16
R9385 VSS.n14526 VSS.n14525 16
R9386 VSS.n14525 VSS.n14524 16
R9387 VSS.n14524 VSS.n14523 16
R9388 VSS.n14523 VSS.n14522 16
R9389 VSS.n14522 VSS.n14521 16
R9390 VSS.n14521 VSS.n14520 16
R9391 VSS.n14520 VSS.n14519 16
R9392 VSS.n14519 VSS.n14518 16
R9393 VSS.n14517 VSS.n14516 16
R9394 VSS.n17091 VSS.n17090 16
R9395 VSS.n17090 VSS.n17089 16
R9396 VSS.n17089 VSS.n17088 16
R9397 VSS.n17088 VSS.n17087 16
R9398 VSS.n17087 VSS.n17086 16
R9399 VSS.n17086 VSS.n17085 16
R9400 VSS.n17085 VSS.n17084 16
R9401 VSS.n17084 VSS.n17083 16
R9402 VSS.n14538 VSS.n14537 16
R9403 VSS.n14537 VSS.n14536 16
R9404 VSS.n14536 VSS.n14535 16
R9405 VSS.n14535 VSS.n14534 16
R9406 VSS.n14534 VSS.n14533 16
R9407 VSS.n14533 VSS.n14532 16
R9408 VSS.n14532 VSS.n14531 16
R9409 VSS.n14531 VSS.n14530 16
R9410 VSS.n14529 VSS.n14528 16
R9411 VSS.n16923 VSS.n16922 16
R9412 VSS.n16922 VSS.n16921 16
R9413 VSS.n16921 VSS.n16920 16
R9414 VSS.n16920 VSS.n16919 16
R9415 VSS.n16919 VSS.n16918 16
R9416 VSS.n16918 VSS.n16917 16
R9417 VSS.n16917 VSS.n16916 16
R9418 VSS.n16916 VSS.n16915 16
R9419 VSS.n14550 VSS.n14549 16
R9420 VSS.n14549 VSS.n14548 16
R9421 VSS.n14548 VSS.n14547 16
R9422 VSS.n14547 VSS.n14546 16
R9423 VSS.n14546 VSS.n14545 16
R9424 VSS.n14545 VSS.n14544 16
R9425 VSS.n14544 VSS.n14543 16
R9426 VSS.n14543 VSS.n14542 16
R9427 VSS.n14541 VSS.n14540 16
R9428 VSS.n16755 VSS.n16754 16
R9429 VSS.n16754 VSS.n16753 16
R9430 VSS.n16753 VSS.n16752 16
R9431 VSS.n16752 VSS.n16751 16
R9432 VSS.n16751 VSS.n16750 16
R9433 VSS.n16750 VSS.n16749 16
R9434 VSS.n16749 VSS.n16748 16
R9435 VSS.n16748 VSS.n16747 16
R9436 VSS.n14075 VSS.n14073 16
R9437 VSS.n14073 VSS.n14072 16
R9438 VSS.n14072 VSS.n14071 16
R9439 VSS.n14071 VSS.n14070 16
R9440 VSS.n14070 VSS.n14069 16
R9441 VSS.n14069 VSS.n14068 16
R9442 VSS.n14068 VSS.n14067 16
R9443 VSS.n14067 VSS.n14066 16
R9444 VSS.n14065 VSS.n14064 16
R9445 VSS.n13907 VSS.n13905 16
R9446 VSS.n13905 VSS.n13904 16
R9447 VSS.n13904 VSS.n13903 16
R9448 VSS.n13903 VSS.n13902 16
R9449 VSS.n13902 VSS.n13901 16
R9450 VSS.n13901 VSS.n13900 16
R9451 VSS.n13900 VSS.n13899 16
R9452 VSS.n13899 VSS.n13898 16
R9453 VSS.n13894 VSS.n13892 16
R9454 VSS.n13892 VSS.n13891 16
R9455 VSS.n13891 VSS.n13890 16
R9456 VSS.n13890 VSS.n13889 16
R9457 VSS.n13889 VSS.n13888 16
R9458 VSS.n13888 VSS.n13887 16
R9459 VSS.n13887 VSS.n13886 16
R9460 VSS.n13886 VSS.n13885 16
R9461 VSS.n13884 VSS.n13883 16
R9462 VSS.n13727 VSS.n13725 16
R9463 VSS.n13725 VSS.n13724 16
R9464 VSS.n13724 VSS.n13723 16
R9465 VSS.n13723 VSS.n13722 16
R9466 VSS.n13722 VSS.n13721 16
R9467 VSS.n13721 VSS.n13720 16
R9468 VSS.n13720 VSS.n13719 16
R9469 VSS.n13719 VSS.n13718 16
R9470 VSS.n13714 VSS.n13712 16
R9471 VSS.n13712 VSS.n13711 16
R9472 VSS.n13711 VSS.n13710 16
R9473 VSS.n13710 VSS.n13709 16
R9474 VSS.n13709 VSS.n13708 16
R9475 VSS.n13708 VSS.n13707 16
R9476 VSS.n13707 VSS.n13706 16
R9477 VSS.n13706 VSS.n13705 16
R9478 VSS.n13704 VSS.n13703 16
R9479 VSS.n13547 VSS.n13545 16
R9480 VSS.n13545 VSS.n13544 16
R9481 VSS.n13544 VSS.n13543 16
R9482 VSS.n13543 VSS.n13542 16
R9483 VSS.n13542 VSS.n13541 16
R9484 VSS.n13541 VSS.n13540 16
R9485 VSS.n13540 VSS.n13539 16
R9486 VSS.n13539 VSS.n13538 16
R9487 VSS.n13534 VSS.n13532 16
R9488 VSS.n13532 VSS.n13531 16
R9489 VSS.n13531 VSS.n13530 16
R9490 VSS.n13530 VSS.n13529 16
R9491 VSS.n13529 VSS.n13528 16
R9492 VSS.n13528 VSS.n13527 16
R9493 VSS.n13527 VSS.n13526 16
R9494 VSS.n13526 VSS.n13525 16
R9495 VSS.n13524 VSS.n13523 16
R9496 VSS.n13367 VSS.n13365 16
R9497 VSS.n13365 VSS.n13364 16
R9498 VSS.n13364 VSS.n13363 16
R9499 VSS.n13363 VSS.n13362 16
R9500 VSS.n13362 VSS.n13361 16
R9501 VSS.n13361 VSS.n13360 16
R9502 VSS.n13360 VSS.n13359 16
R9503 VSS.n13359 VSS.n13358 16
R9504 VSS.n13354 VSS.n13352 16
R9505 VSS.n13352 VSS.n13351 16
R9506 VSS.n13351 VSS.n13350 16
R9507 VSS.n13350 VSS.n13349 16
R9508 VSS.n13349 VSS.n13348 16
R9509 VSS.n13348 VSS.n13347 16
R9510 VSS.n13347 VSS.n13346 16
R9511 VSS.n13346 VSS.n13345 16
R9512 VSS.n13344 VSS.n13343 16
R9513 VSS.n13187 VSS.n13185 16
R9514 VSS.n13185 VSS.n13184 16
R9515 VSS.n13184 VSS.n13183 16
R9516 VSS.n13183 VSS.n13182 16
R9517 VSS.n13182 VSS.n13181 16
R9518 VSS.n13181 VSS.n13180 16
R9519 VSS.n13180 VSS.n13179 16
R9520 VSS.n13179 VSS.n13178 16
R9521 VSS.n13174 VSS.n13172 16
R9522 VSS.n13172 VSS.n13171 16
R9523 VSS.n13171 VSS.n13170 16
R9524 VSS.n13170 VSS.n13169 16
R9525 VSS.n13169 VSS.n13168 16
R9526 VSS.n13168 VSS.n13167 16
R9527 VSS.n13167 VSS.n13166 16
R9528 VSS.n13166 VSS.n13165 16
R9529 VSS.n13164 VSS.n13163 16
R9530 VSS.n13007 VSS.n13005 16
R9531 VSS.n13005 VSS.n13004 16
R9532 VSS.n13004 VSS.n13003 16
R9533 VSS.n13003 VSS.n13002 16
R9534 VSS.n13002 VSS.n13001 16
R9535 VSS.n13001 VSS.n13000 16
R9536 VSS.n13000 VSS.n12999 16
R9537 VSS.n12999 VSS.n12998 16
R9538 VSS.n12994 VSS.n12992 16
R9539 VSS.n12992 VSS.n12991 16
R9540 VSS.n12991 VSS.n12990 16
R9541 VSS.n12990 VSS.n12989 16
R9542 VSS.n12989 VSS.n12988 16
R9543 VSS.n12988 VSS.n12987 16
R9544 VSS.n12987 VSS.n12986 16
R9545 VSS.n12986 VSS.n12985 16
R9546 VSS.n12984 VSS.n12983 16
R9547 VSS.n12827 VSS.n12825 16
R9548 VSS.n12825 VSS.n12824 16
R9549 VSS.n12824 VSS.n12823 16
R9550 VSS.n12823 VSS.n12822 16
R9551 VSS.n12822 VSS.n12821 16
R9552 VSS.n12821 VSS.n12820 16
R9553 VSS.n12820 VSS.n12819 16
R9554 VSS.n12819 VSS.n12818 16
R9555 VSS.n12814 VSS.n12812 16
R9556 VSS.n12812 VSS.n12811 16
R9557 VSS.n12811 VSS.n12810 16
R9558 VSS.n12810 VSS.n12809 16
R9559 VSS.n12809 VSS.n12808 16
R9560 VSS.n12808 VSS.n12807 16
R9561 VSS.n12807 VSS.n12806 16
R9562 VSS.n12806 VSS.n12805 16
R9563 VSS.n12804 VSS.n12803 16
R9564 VSS.n12648 VSS.n12646 16
R9565 VSS.n12646 VSS.n12645 16
R9566 VSS.n12645 VSS.n12644 16
R9567 VSS.n12644 VSS.n12643 16
R9568 VSS.n12643 VSS.n12642 16
R9569 VSS.n12642 VSS.n12641 16
R9570 VSS.n12641 VSS.n12640 16
R9571 VSS.n12640 VSS.n12639 16
R9572 VSS.n9218 VSS.n9216 16
R9573 VSS.n9216 VSS.n9215 16
R9574 VSS.n9215 VSS.n9214 16
R9575 VSS.n9214 VSS.n9213 16
R9576 VSS.n9213 VSS.n9212 16
R9577 VSS.n9212 VSS.n9211 16
R9578 VSS.n9211 VSS.n9210 16
R9579 VSS.n9210 VSS.n9209 16
R9580 VSS.n9208 VSS.n9207 16
R9581 VSS.n7167 VSS.n7165 16
R9582 VSS.n7165 VSS.n7164 16
R9583 VSS.n7164 VSS.n7163 16
R9584 VSS.n7163 VSS.n7162 16
R9585 VSS.n7162 VSS.n7161 16
R9586 VSS.n7161 VSS.n7160 16
R9587 VSS.n7160 VSS.n7159 16
R9588 VSS.n7159 VSS.n7158 16
R9589 VSS.n9386 VSS.n9384 16
R9590 VSS.n9384 VSS.n9383 16
R9591 VSS.n9383 VSS.n9382 16
R9592 VSS.n9382 VSS.n9381 16
R9593 VSS.n9381 VSS.n9380 16
R9594 VSS.n9380 VSS.n9379 16
R9595 VSS.n9379 VSS.n9378 16
R9596 VSS.n9378 VSS.n9377 16
R9597 VSS.n9376 VSS.n9375 16
R9598 VSS.n7155 VSS.n7153 16
R9599 VSS.n7153 VSS.n7152 16
R9600 VSS.n7152 VSS.n7151 16
R9601 VSS.n7151 VSS.n7150 16
R9602 VSS.n7150 VSS.n7149 16
R9603 VSS.n7149 VSS.n7148 16
R9604 VSS.n7148 VSS.n7147 16
R9605 VSS.n7147 VSS.n7146 16
R9606 VSS.n9554 VSS.n9552 16
R9607 VSS.n9552 VSS.n9551 16
R9608 VSS.n9551 VSS.n9550 16
R9609 VSS.n9550 VSS.n9549 16
R9610 VSS.n9549 VSS.n9548 16
R9611 VSS.n9548 VSS.n9547 16
R9612 VSS.n9547 VSS.n9546 16
R9613 VSS.n9546 VSS.n9545 16
R9614 VSS.n9544 VSS.n9543 16
R9615 VSS.n7143 VSS.n7141 16
R9616 VSS.n7141 VSS.n7140 16
R9617 VSS.n7140 VSS.n7139 16
R9618 VSS.n7139 VSS.n7138 16
R9619 VSS.n7138 VSS.n7137 16
R9620 VSS.n7137 VSS.n7136 16
R9621 VSS.n7136 VSS.n7135 16
R9622 VSS.n7135 VSS.n7134 16
R9623 VSS.n9722 VSS.n9720 16
R9624 VSS.n9720 VSS.n9719 16
R9625 VSS.n9719 VSS.n9718 16
R9626 VSS.n9718 VSS.n9717 16
R9627 VSS.n9717 VSS.n9716 16
R9628 VSS.n9716 VSS.n9715 16
R9629 VSS.n9715 VSS.n9714 16
R9630 VSS.n9714 VSS.n9713 16
R9631 VSS.n9712 VSS.n9711 16
R9632 VSS.n7131 VSS.n7129 16
R9633 VSS.n7129 VSS.n7128 16
R9634 VSS.n7128 VSS.n7127 16
R9635 VSS.n7127 VSS.n7126 16
R9636 VSS.n7126 VSS.n7125 16
R9637 VSS.n7125 VSS.n7124 16
R9638 VSS.n7124 VSS.n7123 16
R9639 VSS.n7123 VSS.n7122 16
R9640 VSS.n9890 VSS.n9888 16
R9641 VSS.n9888 VSS.n9887 16
R9642 VSS.n9887 VSS.n9886 16
R9643 VSS.n9886 VSS.n9885 16
R9644 VSS.n9885 VSS.n9884 16
R9645 VSS.n9884 VSS.n9883 16
R9646 VSS.n9883 VSS.n9882 16
R9647 VSS.n9882 VSS.n9881 16
R9648 VSS.n9880 VSS.n9879 16
R9649 VSS.n7119 VSS.n7117 16
R9650 VSS.n7117 VSS.n7116 16
R9651 VSS.n7116 VSS.n7115 16
R9652 VSS.n7115 VSS.n7114 16
R9653 VSS.n7114 VSS.n7113 16
R9654 VSS.n7113 VSS.n7112 16
R9655 VSS.n7112 VSS.n7111 16
R9656 VSS.n7111 VSS.n7110 16
R9657 VSS.n10058 VSS.n10056 16
R9658 VSS.n10056 VSS.n10055 16
R9659 VSS.n10055 VSS.n10054 16
R9660 VSS.n10054 VSS.n10053 16
R9661 VSS.n10053 VSS.n10052 16
R9662 VSS.n10052 VSS.n10051 16
R9663 VSS.n10051 VSS.n10050 16
R9664 VSS.n10050 VSS.n10049 16
R9665 VSS.n10048 VSS.n10047 16
R9666 VSS.n7107 VSS.n7105 16
R9667 VSS.n7105 VSS.n7104 16
R9668 VSS.n7104 VSS.n7103 16
R9669 VSS.n7103 VSS.n7102 16
R9670 VSS.n7102 VSS.n7101 16
R9671 VSS.n7101 VSS.n7100 16
R9672 VSS.n7100 VSS.n7099 16
R9673 VSS.n7099 VSS.n7098 16
R9674 VSS.n10226 VSS.n10224 16
R9675 VSS.n10224 VSS.n10223 16
R9676 VSS.n10223 VSS.n10222 16
R9677 VSS.n10222 VSS.n10221 16
R9678 VSS.n10221 VSS.n10220 16
R9679 VSS.n10220 VSS.n10219 16
R9680 VSS.n10219 VSS.n10218 16
R9681 VSS.n10218 VSS.n10217 16
R9682 VSS.n10216 VSS.n10215 16
R9683 VSS.n7095 VSS.n7093 16
R9684 VSS.n7093 VSS.n7092 16
R9685 VSS.n7092 VSS.n7091 16
R9686 VSS.n7091 VSS.n7090 16
R9687 VSS.n7090 VSS.n7089 16
R9688 VSS.n7089 VSS.n7088 16
R9689 VSS.n7088 VSS.n7087 16
R9690 VSS.n7087 VSS.n7086 16
R9691 VSS.n10393 VSS.n10392 16
R9692 VSS.n10392 VSS.n10391 16
R9693 VSS.n10391 VSS.n10390 16
R9694 VSS.n10390 VSS.n10389 16
R9695 VSS.n10389 VSS.n10388 16
R9696 VSS.n10388 VSS.n10387 16
R9697 VSS.n10387 VSS.n10386 16
R9698 VSS.n10386 VSS.n10385 16
R9699 VSS.n10552 VSS.n10551 16
R9700 VSS.n10384 VSS.n10383 16
R9701 VSS.n10561 VSS.n10560 16
R9702 VSS.n10560 VSS.n10559 16
R9703 VSS.n10559 VSS.n10558 16
R9704 VSS.n10558 VSS.n10557 16
R9705 VSS.n10557 VSS.n10556 16
R9706 VSS.n10556 VSS.n10555 16
R9707 VSS.n10555 VSS.n10554 16
R9708 VSS.n10554 VSS.n10553 16
R9709 VSS.n2461 VSS.n2287 16
R9710 VSS.n2327 VSS.n2287 16
R9711 VSS.n2330 VSS.n2327 16
R9712 VSS.n2331 VSS.n2330 16
R9713 VSS.n2334 VSS.n2331 16
R9714 VSS.n2335 VSS.n2334 16
R9715 VSS.n2338 VSS.n2335 16
R9716 VSS.n2340 VSS.n2338 16
R9717 VSS.n2356 VSS.n2355 16
R9718 VSS.n2355 VSS.n2352 16
R9719 VSS.n2352 VSS.n2351 16
R9720 VSS.n2351 VSS.n2348 16
R9721 VSS.n2348 VSS.n2347 16
R9722 VSS.n2347 VSS.n2344 16
R9723 VSS.n2344 VSS.n2343 16
R9724 VSS.n2343 VSS.n2341 16
R9725 VSS.n2374 VSS.n2373 16
R9726 VSS.n2373 VSS.n2371 16
R9727 VSS.n2371 VSS.n2368 16
R9728 VSS.n2368 VSS.n2367 16
R9729 VSS.n2367 VSS.n2364 16
R9730 VSS.n2364 VSS.n2363 16
R9731 VSS.n2363 VSS.n2360 16
R9732 VSS.n2360 VSS.n2359 16
R9733 VSS.n2551 VSS.n2197 16
R9734 VSS.n2237 VSS.n2197 16
R9735 VSS.n2240 VSS.n2237 16
R9736 VSS.n2241 VSS.n2240 16
R9737 VSS.n2244 VSS.n2241 16
R9738 VSS.n2245 VSS.n2244 16
R9739 VSS.n2248 VSS.n2245 16
R9740 VSS.n2250 VSS.n2248 16
R9741 VSS.n2266 VSS.n2265 16
R9742 VSS.n2265 VSS.n2262 16
R9743 VSS.n2262 VSS.n2261 16
R9744 VSS.n2261 VSS.n2258 16
R9745 VSS.n2258 VSS.n2257 16
R9746 VSS.n2257 VSS.n2254 16
R9747 VSS.n2254 VSS.n2253 16
R9748 VSS.n2253 VSS.n2251 16
R9749 VSS.n2284 VSS.n2283 16
R9750 VSS.n2283 VSS.n2281 16
R9751 VSS.n2281 VSS.n2278 16
R9752 VSS.n2278 VSS.n2277 16
R9753 VSS.n2277 VSS.n2274 16
R9754 VSS.n2274 VSS.n2273 16
R9755 VSS.n2273 VSS.n2270 16
R9756 VSS.n2270 VSS.n2269 16
R9757 VSS.n2641 VSS.n2107 16
R9758 VSS.n2147 VSS.n2107 16
R9759 VSS.n2150 VSS.n2147 16
R9760 VSS.n2151 VSS.n2150 16
R9761 VSS.n2154 VSS.n2151 16
R9762 VSS.n2155 VSS.n2154 16
R9763 VSS.n2158 VSS.n2155 16
R9764 VSS.n2160 VSS.n2158 16
R9765 VSS.n2176 VSS.n2175 16
R9766 VSS.n2175 VSS.n2172 16
R9767 VSS.n2172 VSS.n2171 16
R9768 VSS.n2171 VSS.n2168 16
R9769 VSS.n2168 VSS.n2167 16
R9770 VSS.n2167 VSS.n2164 16
R9771 VSS.n2164 VSS.n2163 16
R9772 VSS.n2163 VSS.n2161 16
R9773 VSS.n2194 VSS.n2193 16
R9774 VSS.n2193 VSS.n2191 16
R9775 VSS.n2191 VSS.n2188 16
R9776 VSS.n2188 VSS.n2187 16
R9777 VSS.n2187 VSS.n2184 16
R9778 VSS.n2184 VSS.n2183 16
R9779 VSS.n2183 VSS.n2180 16
R9780 VSS.n2180 VSS.n2179 16
R9781 VSS.n2731 VSS.n2017 16
R9782 VSS.n2057 VSS.n2017 16
R9783 VSS.n2060 VSS.n2057 16
R9784 VSS.n2061 VSS.n2060 16
R9785 VSS.n2064 VSS.n2061 16
R9786 VSS.n2065 VSS.n2064 16
R9787 VSS.n2068 VSS.n2065 16
R9788 VSS.n2070 VSS.n2068 16
R9789 VSS.n2086 VSS.n2085 16
R9790 VSS.n2085 VSS.n2082 16
R9791 VSS.n2082 VSS.n2081 16
R9792 VSS.n2081 VSS.n2078 16
R9793 VSS.n2078 VSS.n2077 16
R9794 VSS.n2077 VSS.n2074 16
R9795 VSS.n2074 VSS.n2073 16
R9796 VSS.n2073 VSS.n2071 16
R9797 VSS.n2104 VSS.n2103 16
R9798 VSS.n2103 VSS.n2101 16
R9799 VSS.n2101 VSS.n2098 16
R9800 VSS.n2098 VSS.n2097 16
R9801 VSS.n2097 VSS.n2094 16
R9802 VSS.n2094 VSS.n2093 16
R9803 VSS.n2093 VSS.n2090 16
R9804 VSS.n2090 VSS.n2089 16
R9805 VSS.n2821 VSS.n1927 16
R9806 VSS.n1967 VSS.n1927 16
R9807 VSS.n1970 VSS.n1967 16
R9808 VSS.n1971 VSS.n1970 16
R9809 VSS.n1974 VSS.n1971 16
R9810 VSS.n1975 VSS.n1974 16
R9811 VSS.n1978 VSS.n1975 16
R9812 VSS.n1980 VSS.n1978 16
R9813 VSS.n1996 VSS.n1995 16
R9814 VSS.n1995 VSS.n1992 16
R9815 VSS.n1992 VSS.n1991 16
R9816 VSS.n1991 VSS.n1988 16
R9817 VSS.n1988 VSS.n1987 16
R9818 VSS.n1987 VSS.n1984 16
R9819 VSS.n1984 VSS.n1983 16
R9820 VSS.n1983 VSS.n1981 16
R9821 VSS.n2014 VSS.n2013 16
R9822 VSS.n2013 VSS.n2011 16
R9823 VSS.n2011 VSS.n2008 16
R9824 VSS.n2008 VSS.n2007 16
R9825 VSS.n2007 VSS.n2004 16
R9826 VSS.n2004 VSS.n2003 16
R9827 VSS.n2003 VSS.n2000 16
R9828 VSS.n2000 VSS.n1999 16
R9829 VSS.n2911 VSS.n1837 16
R9830 VSS.n1877 VSS.n1837 16
R9831 VSS.n1880 VSS.n1877 16
R9832 VSS.n1881 VSS.n1880 16
R9833 VSS.n1884 VSS.n1881 16
R9834 VSS.n1885 VSS.n1884 16
R9835 VSS.n1888 VSS.n1885 16
R9836 VSS.n1890 VSS.n1888 16
R9837 VSS.n1906 VSS.n1905 16
R9838 VSS.n1905 VSS.n1902 16
R9839 VSS.n1902 VSS.n1901 16
R9840 VSS.n1901 VSS.n1898 16
R9841 VSS.n1898 VSS.n1897 16
R9842 VSS.n1897 VSS.n1894 16
R9843 VSS.n1894 VSS.n1893 16
R9844 VSS.n1893 VSS.n1891 16
R9845 VSS.n1924 VSS.n1923 16
R9846 VSS.n1923 VSS.n1921 16
R9847 VSS.n1921 VSS.n1918 16
R9848 VSS.n1918 VSS.n1917 16
R9849 VSS.n1917 VSS.n1914 16
R9850 VSS.n1914 VSS.n1913 16
R9851 VSS.n1913 VSS.n1910 16
R9852 VSS.n1910 VSS.n1909 16
R9853 VSS.n3001 VSS.n1747 16
R9854 VSS.n1787 VSS.n1747 16
R9855 VSS.n1790 VSS.n1787 16
R9856 VSS.n1791 VSS.n1790 16
R9857 VSS.n1794 VSS.n1791 16
R9858 VSS.n1795 VSS.n1794 16
R9859 VSS.n1798 VSS.n1795 16
R9860 VSS.n1800 VSS.n1798 16
R9861 VSS.n1816 VSS.n1815 16
R9862 VSS.n1815 VSS.n1812 16
R9863 VSS.n1812 VSS.n1811 16
R9864 VSS.n1811 VSS.n1808 16
R9865 VSS.n1808 VSS.n1807 16
R9866 VSS.n1807 VSS.n1804 16
R9867 VSS.n1804 VSS.n1803 16
R9868 VSS.n1803 VSS.n1801 16
R9869 VSS.n1834 VSS.n1833 16
R9870 VSS.n1833 VSS.n1831 16
R9871 VSS.n1831 VSS.n1828 16
R9872 VSS.n1828 VSS.n1827 16
R9873 VSS.n1827 VSS.n1824 16
R9874 VSS.n1824 VSS.n1823 16
R9875 VSS.n1823 VSS.n1820 16
R9876 VSS.n1820 VSS.n1819 16
R9877 VSS.n3091 VSS.n1657 16
R9878 VSS.n1697 VSS.n1657 16
R9879 VSS.n1700 VSS.n1697 16
R9880 VSS.n1701 VSS.n1700 16
R9881 VSS.n1704 VSS.n1701 16
R9882 VSS.n1705 VSS.n1704 16
R9883 VSS.n1708 VSS.n1705 16
R9884 VSS.n1710 VSS.n1708 16
R9885 VSS.n1726 VSS.n1725 16
R9886 VSS.n1725 VSS.n1722 16
R9887 VSS.n1722 VSS.n1721 16
R9888 VSS.n1721 VSS.n1718 16
R9889 VSS.n1718 VSS.n1717 16
R9890 VSS.n1717 VSS.n1714 16
R9891 VSS.n1714 VSS.n1713 16
R9892 VSS.n1713 VSS.n1711 16
R9893 VSS.n1744 VSS.n1743 16
R9894 VSS.n1743 VSS.n1741 16
R9895 VSS.n1741 VSS.n1738 16
R9896 VSS.n1738 VSS.n1737 16
R9897 VSS.n1737 VSS.n1734 16
R9898 VSS.n1734 VSS.n1733 16
R9899 VSS.n1733 VSS.n1730 16
R9900 VSS.n1730 VSS.n1729 16
R9901 VSS.n6239 VSS.n6238 16
R9902 VSS.n6238 VSS.n6235 16
R9903 VSS.n6235 VSS.n6234 16
R9904 VSS.n6234 VSS.n6231 16
R9905 VSS.n6231 VSS.n6230 16
R9906 VSS.n6230 VSS.n6227 16
R9907 VSS.n6227 VSS.n6226 16
R9908 VSS.n6226 VSS.n6223 16
R9909 VSS.n6207 VSS.n6206 16
R9910 VSS.n6210 VSS.n6207 16
R9911 VSS.n6211 VSS.n6210 16
R9912 VSS.n6214 VSS.n6211 16
R9913 VSS.n6215 VSS.n6214 16
R9914 VSS.n6218 VSS.n6215 16
R9915 VSS.n6219 VSS.n6218 16
R9916 VSS.n6222 VSS.n6219 16
R9917 VSS.n6190 VSS.n6074 16
R9918 VSS.n6193 VSS.n6190 16
R9919 VSS.n6194 VSS.n6193 16
R9920 VSS.n6197 VSS.n6194 16
R9921 VSS.n6198 VSS.n6197 16
R9922 VSS.n6201 VSS.n6198 16
R9923 VSS.n6203 VSS.n6201 16
R9924 VSS.n6204 VSS.n6203 16
R9925 VSS.n6303 VSS.n6302 16
R9926 VSS.n6302 VSS.n6299 16
R9927 VSS.n6299 VSS.n6298 16
R9928 VSS.n6298 VSS.n6295 16
R9929 VSS.n6295 VSS.n6294 16
R9930 VSS.n6294 VSS.n6291 16
R9931 VSS.n6291 VSS.n6290 16
R9932 VSS.n6290 VSS.n6287 16
R9933 VSS.n6271 VSS.n6270 16
R9934 VSS.n6274 VSS.n6271 16
R9935 VSS.n6275 VSS.n6274 16
R9936 VSS.n6278 VSS.n6275 16
R9937 VSS.n6279 VSS.n6278 16
R9938 VSS.n6282 VSS.n6279 16
R9939 VSS.n6283 VSS.n6282 16
R9940 VSS.n6286 VSS.n6283 16
R9941 VSS.n6254 VSS.n5958 16
R9942 VSS.n6257 VSS.n6254 16
R9943 VSS.n6258 VSS.n6257 16
R9944 VSS.n6261 VSS.n6258 16
R9945 VSS.n6262 VSS.n6261 16
R9946 VSS.n6265 VSS.n6262 16
R9947 VSS.n6267 VSS.n6265 16
R9948 VSS.n6268 VSS.n6267 16
R9949 VSS.n6367 VSS.n6366 16
R9950 VSS.n6366 VSS.n6363 16
R9951 VSS.n6363 VSS.n6362 16
R9952 VSS.n6362 VSS.n6359 16
R9953 VSS.n6359 VSS.n6358 16
R9954 VSS.n6358 VSS.n6355 16
R9955 VSS.n6355 VSS.n6354 16
R9956 VSS.n6354 VSS.n6351 16
R9957 VSS.n6335 VSS.n6334 16
R9958 VSS.n6338 VSS.n6335 16
R9959 VSS.n6339 VSS.n6338 16
R9960 VSS.n6342 VSS.n6339 16
R9961 VSS.n6343 VSS.n6342 16
R9962 VSS.n6346 VSS.n6343 16
R9963 VSS.n6347 VSS.n6346 16
R9964 VSS.n6350 VSS.n6347 16
R9965 VSS.n6318 VSS.n5842 16
R9966 VSS.n6321 VSS.n6318 16
R9967 VSS.n6322 VSS.n6321 16
R9968 VSS.n6325 VSS.n6322 16
R9969 VSS.n6326 VSS.n6325 16
R9970 VSS.n6329 VSS.n6326 16
R9971 VSS.n6331 VSS.n6329 16
R9972 VSS.n6332 VSS.n6331 16
R9973 VSS.n6990 VSS.n6383 16
R9974 VSS.n6990 VSS.n6989 16
R9975 VSS.n6989 VSS.n6988 16
R9976 VSS.n6988 VSS.n6385 16
R9977 VSS.n6983 VSS.n6385 16
R9978 VSS.n6983 VSS.n6982 16
R9979 VSS.n6982 VSS.n6981 16
R9980 VSS.n6981 VSS.n6388 16
R9981 VSS.n6960 VSS.n6393 16
R9982 VSS.n6966 VSS.n6393 16
R9983 VSS.n6967 VSS.n6966 16
R9984 VSS.n6968 VSS.n6967 16
R9985 VSS.n6968 VSS.n6391 16
R9986 VSS.n6974 VSS.n6391 16
R9987 VSS.n6975 VSS.n6974 16
R9988 VSS.n6976 VSS.n6975 16
R9989 VSS.n6946 VSS.n6945 16
R9990 VSS.n6947 VSS.n6946 16
R9991 VSS.n6947 VSS.n6397 16
R9992 VSS.n6952 VSS.n6397 16
R9993 VSS.n6953 VSS.n6952 16
R9994 VSS.n6953 VSS.n6395 16
R9995 VSS.n6958 VSS.n6395 16
R9996 VSS.n6959 VSS.n6958 16
R9997 VSS.n6935 VSS.n6401 16
R9998 VSS.n6441 VSS.n6401 16
R9999 VSS.n6444 VSS.n6441 16
R10000 VSS.n6445 VSS.n6444 16
R10001 VSS.n6448 VSS.n6445 16
R10002 VSS.n6449 VSS.n6448 16
R10003 VSS.n6452 VSS.n6449 16
R10004 VSS.n6454 VSS.n6452 16
R10005 VSS.n6470 VSS.n6469 16
R10006 VSS.n6469 VSS.n6466 16
R10007 VSS.n6466 VSS.n6465 16
R10008 VSS.n6465 VSS.n6462 16
R10009 VSS.n6462 VSS.n6461 16
R10010 VSS.n6461 VSS.n6458 16
R10011 VSS.n6458 VSS.n6457 16
R10012 VSS.n6457 VSS.n6455 16
R10013 VSS.n6488 VSS.n6487 16
R10014 VSS.n6487 VSS.n6485 16
R10015 VSS.n6485 VSS.n6482 16
R10016 VSS.n6482 VSS.n6481 16
R10017 VSS.n6481 VSS.n6478 16
R10018 VSS.n6478 VSS.n6477 16
R10019 VSS.n6477 VSS.n6474 16
R10020 VSS.n6474 VSS.n6473 16
R10021 VSS.n6845 VSS.n6491 16
R10022 VSS.n6531 VSS.n6491 16
R10023 VSS.n6534 VSS.n6531 16
R10024 VSS.n6535 VSS.n6534 16
R10025 VSS.n6538 VSS.n6535 16
R10026 VSS.n6539 VSS.n6538 16
R10027 VSS.n6542 VSS.n6539 16
R10028 VSS.n6544 VSS.n6542 16
R10029 VSS.n6560 VSS.n6559 16
R10030 VSS.n6559 VSS.n6556 16
R10031 VSS.n6556 VSS.n6555 16
R10032 VSS.n6555 VSS.n6552 16
R10033 VSS.n6552 VSS.n6551 16
R10034 VSS.n6551 VSS.n6548 16
R10035 VSS.n6548 VSS.n6547 16
R10036 VSS.n6547 VSS.n6545 16
R10037 VSS.n6578 VSS.n6577 16
R10038 VSS.n6577 VSS.n6575 16
R10039 VSS.n6575 VSS.n6572 16
R10040 VSS.n6572 VSS.n6571 16
R10041 VSS.n6571 VSS.n6568 16
R10042 VSS.n6568 VSS.n6567 16
R10043 VSS.n6567 VSS.n6564 16
R10044 VSS.n6564 VSS.n6563 16
R10045 VSS.n6755 VSS.n6581 16
R10046 VSS.n6621 VSS.n6581 16
R10047 VSS.n6624 VSS.n6621 16
R10048 VSS.n6625 VSS.n6624 16
R10049 VSS.n6628 VSS.n6625 16
R10050 VSS.n6629 VSS.n6628 16
R10051 VSS.n6632 VSS.n6629 16
R10052 VSS.n6634 VSS.n6632 16
R10053 VSS.n6650 VSS.n6649 16
R10054 VSS.n6649 VSS.n6646 16
R10055 VSS.n6646 VSS.n6645 16
R10056 VSS.n6645 VSS.n6642 16
R10057 VSS.n6642 VSS.n6641 16
R10058 VSS.n6641 VSS.n6638 16
R10059 VSS.n6638 VSS.n6637 16
R10060 VSS.n6637 VSS.n6635 16
R10061 VSS.n6668 VSS.n6667 16
R10062 VSS.n6667 VSS.n6665 16
R10063 VSS.n6665 VSS.n6662 16
R10064 VSS.n6662 VSS.n6661 16
R10065 VSS.n6661 VSS.n6658 16
R10066 VSS.n6658 VSS.n6657 16
R10067 VSS.n6657 VSS.n6654 16
R10068 VSS.n6654 VSS.n6653 16
R10069 VSS.n18000 VSS.n17998 16
R10070 VSS.n18002 VSS.n18000 16
R10071 VSS.n18004 VSS.n18002 16
R10072 VSS.n18006 VSS.n18004 16
R10073 VSS.n18008 VSS.n18006 16
R10074 VSS.n18010 VSS.n18008 16
R10075 VSS.n18012 VSS.n18010 16
R10076 VSS.n18013 VSS.n18012 16
R10077 VSS.n17996 VSS.n17993 16
R10078 VSS.n17993 VSS.n17992 16
R10079 VSS.n17992 VSS.n17989 16
R10080 VSS.n17989 VSS.n17988 16
R10081 VSS.n17988 VSS.n17985 16
R10082 VSS.n17984 VSS.n17981 16
R10083 VSS.n17981 VSS.n17980 16
R10084 VSS.n17977 VSS.n17976 16
R10085 VSS.n17976 VSS.n17973 16
R10086 VSS.n17973 VSS.n17972 16
R10087 VSS.n17972 VSS.n17969 16
R10088 VSS.n17969 VSS.n17968 16
R10089 VSS.n17968 VSS.n17965 16
R10090 VSS.n17965 VSS.n17964 16
R10091 VSS.n17964 VSS.n17961 16
R10092 VSS.n18014 VSS.n17922 16
R10093 VSS.n17952 VSS.n17949 16
R10094 VSS.n17953 VSS.n17952 16
R10095 VSS.n17956 VSS.n17953 16
R10096 VSS.n17957 VSS.n17956 16
R10097 VSS.n17960 VSS.n17957 16
R10098 VSS VSS.n7058 15.813
R10099 VSS.n14096 VSS.n14095 15.375
R10100 VSS.n2462 VSS.n2286 14.755
R10101 VSS.n2552 VSS.n2196 14.755
R10102 VSS.n2642 VSS.n2106 14.755
R10103 VSS.n2732 VSS.n2016 14.755
R10104 VSS.n2822 VSS.n1926 14.755
R10105 VSS.n2912 VSS.n1836 14.755
R10106 VSS.n3002 VSS.n1746 14.755
R10107 VSS.n3092 VSS.n1656 14.755
R10108 VSS.n6241 VSS.n6240 14.755
R10109 VSS.n6305 VSS.n6304 14.755
R10110 VSS.n6369 VSS.n6368 14.755
R10111 VSS.n6382 VSS.n5838 14.755
R10112 VSS.n6936 VSS.n6400 14.755
R10113 VSS.n6846 VSS.n6490 14.755
R10114 VSS.n6756 VSS.n6580 14.755
R10115 VSS.n14459 VSS.n14413 14.615
R10116 VSS.n14279 VSS.n14233 14.615
R10117 VSS.n14056 VSS.n14010 14.615
R10118 VSS.n13876 VSS.n13830 14.615
R10119 VSS.n13696 VSS.n13650 14.615
R10120 VSS.n13516 VSS.n13470 14.615
R10121 VSS.n13336 VSS.n13290 14.615
R10122 VSS.n13156 VSS.n13110 14.615
R10123 VSS.n12976 VSS.n12930 14.615
R10124 VSS.n12796 VSS.n12750 14.615
R10125 VSS.n9226 VSS.n9225 14.615
R10126 VSS.n9394 VSS.n9393 14.615
R10127 VSS.n9562 VSS.n9561 14.615
R10128 VSS.n9730 VSS.n9729 14.615
R10129 VSS.n9898 VSS.n9897 14.615
R10130 VSS.n10066 VSS.n10065 14.615
R10131 VSS.n10234 VSS.n10233 14.615
R10132 VSS.n6931 VSS.n6422 14.615
R10133 VSS.n6841 VSS.n6512 14.615
R10134 VSS.n6751 VSS.n6602 14.615
R10135 VSS.n18020 VSS.n17922 13.949
R10136 VSS.n14651 VSS.n14650 13.653
R10137 VSS.n14665 VSS.n14664 13.653
R10138 VSS.n14679 VSS.n14678 13.653
R10139 VSS.n14693 VSS.n14692 13.653
R10140 VSS.n14707 VSS.n14706 13.653
R10141 VSS.n14721 VSS.n14720 13.653
R10142 VSS.n14725 VSS.n14724 13.653
R10143 VSS.n14743 VSS.n14742 13.653
R10144 VSS.n14757 VSS.n14756 13.653
R10145 VSS.n14771 VSS.n14770 13.653
R10146 VSS.n14785 VSS.n14784 13.653
R10147 VSS.n14799 VSS.n14798 13.653
R10148 VSS.n15151 VSS.n15150 13.653
R10149 VSS.n15165 VSS.n15164 13.653
R10150 VSS.n15179 VSS.n15178 13.653
R10151 VSS.n15193 VSS.n15192 13.653
R10152 VSS.n15207 VSS.n15206 13.653
R10153 VSS.n15221 VSS.n15220 13.653
R10154 VSS.n15225 VSS.n15224 13.653
R10155 VSS.n15243 VSS.n15242 13.653
R10156 VSS.n15257 VSS.n15256 13.653
R10157 VSS.n15271 VSS.n15270 13.653
R10158 VSS.n15285 VSS.n15284 13.653
R10159 VSS.n15299 VSS.n15298 13.653
R10160 VSS.n14907 VSS.n14906 13.653
R10161 VSS.n14921 VSS.n14920 13.653
R10162 VSS.n14935 VSS.n14934 13.653
R10163 VSS.n14949 VSS.n14948 13.653
R10164 VSS.n14963 VSS.n14962 13.653
R10165 VSS.n14977 VSS.n14976 13.653
R10166 VSS.n14981 VSS.n14980 13.653
R10167 VSS.n14999 VSS.n14998 13.653
R10168 VSS.n15013 VSS.n15012 13.653
R10169 VSS.n15027 VSS.n15026 13.653
R10170 VSS.n15041 VSS.n15040 13.653
R10171 VSS.n15055 VSS.n15054 13.653
R10172 VSS.n15639 VSS.n15638 13.653
R10173 VSS.n15653 VSS.n15652 13.653
R10174 VSS.n15667 VSS.n15666 13.653
R10175 VSS.n15681 VSS.n15680 13.653
R10176 VSS.n15695 VSS.n15694 13.653
R10177 VSS.n15709 VSS.n15708 13.653
R10178 VSS.n15713 VSS.n15712 13.653
R10179 VSS.n15731 VSS.n15730 13.653
R10180 VSS.n15745 VSS.n15744 13.653
R10181 VSS.n15759 VSS.n15758 13.653
R10182 VSS.n15773 VSS.n15772 13.653
R10183 VSS.n15787 VSS.n15786 13.653
R10184 VSS.n15395 VSS.n15394 13.653
R10185 VSS.n15409 VSS.n15408 13.653
R10186 VSS.n15423 VSS.n15422 13.653
R10187 VSS.n15437 VSS.n15436 13.653
R10188 VSS.n15451 VSS.n15450 13.653
R10189 VSS.n15465 VSS.n15464 13.653
R10190 VSS.n15469 VSS.n15468 13.653
R10191 VSS.n15487 VSS.n15486 13.653
R10192 VSS.n15501 VSS.n15500 13.653
R10193 VSS.n15515 VSS.n15514 13.653
R10194 VSS.n15529 VSS.n15528 13.653
R10195 VSS.n15543 VSS.n15542 13.653
R10196 VSS.n16127 VSS.n16126 13.653
R10197 VSS.n16141 VSS.n16140 13.653
R10198 VSS.n16155 VSS.n16154 13.653
R10199 VSS.n16169 VSS.n16168 13.653
R10200 VSS.n16183 VSS.n16182 13.653
R10201 VSS.n16197 VSS.n16196 13.653
R10202 VSS.n16201 VSS.n16200 13.653
R10203 VSS.n16219 VSS.n16218 13.653
R10204 VSS.n16233 VSS.n16232 13.653
R10205 VSS.n16247 VSS.n16246 13.653
R10206 VSS.n16261 VSS.n16260 13.653
R10207 VSS.n16275 VSS.n16274 13.653
R10208 VSS.n15883 VSS.n15882 13.653
R10209 VSS.n15897 VSS.n15896 13.653
R10210 VSS.n15911 VSS.n15910 13.653
R10211 VSS.n15925 VSS.n15924 13.653
R10212 VSS.n15939 VSS.n15938 13.653
R10213 VSS.n15953 VSS.n15952 13.653
R10214 VSS.n15957 VSS.n15956 13.653
R10215 VSS.n15975 VSS.n15974 13.653
R10216 VSS.n15989 VSS.n15988 13.653
R10217 VSS.n16003 VSS.n16002 13.653
R10218 VSS.n16017 VSS.n16016 13.653
R10219 VSS.n16031 VSS.n16030 13.653
R10220 VSS.n16383 VSS.n16382 13.653
R10221 VSS.n16397 VSS.n16396 13.653
R10222 VSS.n16411 VSS.n16410 13.653
R10223 VSS.n16425 VSS.n16424 13.653
R10224 VSS.n16439 VSS.n16438 13.653
R10225 VSS.n16453 VSS.n16452 13.653
R10226 VSS.n16457 VSS.n16456 13.653
R10227 VSS.n16475 VSS.n16474 13.653
R10228 VSS.n16489 VSS.n16488 13.653
R10229 VSS.n16503 VSS.n16502 13.653
R10230 VSS.n16517 VSS.n16516 13.653
R10231 VSS.n16576 VSS.n16575 13.653
R10232 VSS.n10700 VSS.n10699 13.653
R10233 VSS.n10714 VSS.n10713 13.653
R10234 VSS.n10728 VSS.n10727 13.653
R10235 VSS.n10742 VSS.n10741 13.653
R10236 VSS.n10756 VSS.n10755 13.653
R10237 VSS.n10770 VSS.n10769 13.653
R10238 VSS.n10774 VSS.n10773 13.653
R10239 VSS.n10792 VSS.n10791 13.653
R10240 VSS.n10806 VSS.n10805 13.653
R10241 VSS.n10820 VSS.n10819 13.653
R10242 VSS.n10834 VSS.n10833 13.653
R10243 VSS.n10848 VSS.n10847 13.653
R10244 VSS.n11200 VSS.n11199 13.653
R10245 VSS.n11214 VSS.n11213 13.653
R10246 VSS.n11228 VSS.n11227 13.653
R10247 VSS.n11242 VSS.n11241 13.653
R10248 VSS.n11256 VSS.n11255 13.653
R10249 VSS.n11270 VSS.n11269 13.653
R10250 VSS.n11274 VSS.n11273 13.653
R10251 VSS.n11292 VSS.n11291 13.653
R10252 VSS.n11306 VSS.n11305 13.653
R10253 VSS.n11320 VSS.n11319 13.653
R10254 VSS.n11334 VSS.n11333 13.653
R10255 VSS.n11348 VSS.n11347 13.653
R10256 VSS.n10956 VSS.n10955 13.653
R10257 VSS.n10970 VSS.n10969 13.653
R10258 VSS.n10984 VSS.n10983 13.653
R10259 VSS.n10998 VSS.n10997 13.653
R10260 VSS.n11012 VSS.n11011 13.653
R10261 VSS.n11026 VSS.n11025 13.653
R10262 VSS.n11030 VSS.n11029 13.653
R10263 VSS.n11048 VSS.n11047 13.653
R10264 VSS.n11062 VSS.n11061 13.653
R10265 VSS.n11076 VSS.n11075 13.653
R10266 VSS.n11090 VSS.n11089 13.653
R10267 VSS.n11104 VSS.n11103 13.653
R10268 VSS.n11688 VSS.n11687 13.653
R10269 VSS.n11702 VSS.n11701 13.653
R10270 VSS.n11716 VSS.n11715 13.653
R10271 VSS.n11730 VSS.n11729 13.653
R10272 VSS.n11744 VSS.n11743 13.653
R10273 VSS.n11758 VSS.n11757 13.653
R10274 VSS.n11762 VSS.n11761 13.653
R10275 VSS.n11780 VSS.n11779 13.653
R10276 VSS.n11794 VSS.n11793 13.653
R10277 VSS.n11808 VSS.n11807 13.653
R10278 VSS.n11822 VSS.n11821 13.653
R10279 VSS.n11836 VSS.n11835 13.653
R10280 VSS.n11444 VSS.n11443 13.653
R10281 VSS.n11458 VSS.n11457 13.653
R10282 VSS.n11472 VSS.n11471 13.653
R10283 VSS.n11486 VSS.n11485 13.653
R10284 VSS.n11500 VSS.n11499 13.653
R10285 VSS.n11514 VSS.n11513 13.653
R10286 VSS.n11518 VSS.n11517 13.653
R10287 VSS.n11536 VSS.n11535 13.653
R10288 VSS.n11550 VSS.n11549 13.653
R10289 VSS.n11564 VSS.n11563 13.653
R10290 VSS.n11578 VSS.n11577 13.653
R10291 VSS.n11592 VSS.n11591 13.653
R10292 VSS.n12176 VSS.n12175 13.653
R10293 VSS.n12190 VSS.n12189 13.653
R10294 VSS.n12204 VSS.n12203 13.653
R10295 VSS.n12218 VSS.n12217 13.653
R10296 VSS.n12232 VSS.n12231 13.653
R10297 VSS.n12246 VSS.n12245 13.653
R10298 VSS.n12250 VSS.n12249 13.653
R10299 VSS.n12268 VSS.n12267 13.653
R10300 VSS.n12282 VSS.n12281 13.653
R10301 VSS.n12296 VSS.n12295 13.653
R10302 VSS.n12310 VSS.n12309 13.653
R10303 VSS.n12324 VSS.n12323 13.653
R10304 VSS.n11932 VSS.n11931 13.653
R10305 VSS.n11946 VSS.n11945 13.653
R10306 VSS.n11960 VSS.n11959 13.653
R10307 VSS.n11974 VSS.n11973 13.653
R10308 VSS.n11988 VSS.n11987 13.653
R10309 VSS.n12002 VSS.n12001 13.653
R10310 VSS.n12006 VSS.n12005 13.653
R10311 VSS.n12024 VSS.n12023 13.653
R10312 VSS.n12038 VSS.n12037 13.653
R10313 VSS.n12052 VSS.n12051 13.653
R10314 VSS.n12066 VSS.n12065 13.653
R10315 VSS.n12080 VSS.n12079 13.653
R10316 VSS.n12432 VSS.n12431 13.653
R10317 VSS.n12446 VSS.n12445 13.653
R10318 VSS.n12460 VSS.n12459 13.653
R10319 VSS.n12474 VSS.n12473 13.653
R10320 VSS.n12488 VSS.n12487 13.653
R10321 VSS.n12502 VSS.n12501 13.653
R10322 VSS.n12506 VSS.n12505 13.653
R10323 VSS.n12524 VSS.n12523 13.653
R10324 VSS.n12538 VSS.n12537 13.653
R10325 VSS.n12552 VSS.n12551 13.653
R10326 VSS.n12566 VSS.n12565 13.653
R10327 VSS.n12625 VSS.n12624 13.653
R10328 VSS.n7268 VSS.n7267 13.653
R10329 VSS.n7282 VSS.n7281 13.653
R10330 VSS.n7296 VSS.n7295 13.653
R10331 VSS.n7310 VSS.n7309 13.653
R10332 VSS.n7324 VSS.n7323 13.653
R10333 VSS.n7338 VSS.n7337 13.653
R10334 VSS.n7342 VSS.n7341 13.653
R10335 VSS.n7360 VSS.n7359 13.653
R10336 VSS.n7374 VSS.n7373 13.653
R10337 VSS.n7388 VSS.n7387 13.653
R10338 VSS.n7402 VSS.n7401 13.653
R10339 VSS.n7416 VSS.n7415 13.653
R10340 VSS.n7768 VSS.n7767 13.653
R10341 VSS.n7782 VSS.n7781 13.653
R10342 VSS.n7796 VSS.n7795 13.653
R10343 VSS.n7810 VSS.n7809 13.653
R10344 VSS.n7824 VSS.n7823 13.653
R10345 VSS.n7838 VSS.n7837 13.653
R10346 VSS.n7842 VSS.n7841 13.653
R10347 VSS.n7860 VSS.n7859 13.653
R10348 VSS.n7874 VSS.n7873 13.653
R10349 VSS.n7888 VSS.n7887 13.653
R10350 VSS.n7902 VSS.n7901 13.653
R10351 VSS.n7916 VSS.n7915 13.653
R10352 VSS.n7524 VSS.n7523 13.653
R10353 VSS.n7538 VSS.n7537 13.653
R10354 VSS.n7552 VSS.n7551 13.653
R10355 VSS.n7566 VSS.n7565 13.653
R10356 VSS.n7580 VSS.n7579 13.653
R10357 VSS.n7594 VSS.n7593 13.653
R10358 VSS.n7598 VSS.n7597 13.653
R10359 VSS.n7616 VSS.n7615 13.653
R10360 VSS.n7630 VSS.n7629 13.653
R10361 VSS.n7644 VSS.n7643 13.653
R10362 VSS.n7658 VSS.n7657 13.653
R10363 VSS.n7672 VSS.n7671 13.653
R10364 VSS.n8256 VSS.n8255 13.653
R10365 VSS.n8270 VSS.n8269 13.653
R10366 VSS.n8284 VSS.n8283 13.653
R10367 VSS.n8298 VSS.n8297 13.653
R10368 VSS.n8312 VSS.n8311 13.653
R10369 VSS.n8326 VSS.n8325 13.653
R10370 VSS.n8330 VSS.n8329 13.653
R10371 VSS.n8348 VSS.n8347 13.653
R10372 VSS.n8362 VSS.n8361 13.653
R10373 VSS.n8376 VSS.n8375 13.653
R10374 VSS.n8390 VSS.n8389 13.653
R10375 VSS.n8404 VSS.n8403 13.653
R10376 VSS.n8012 VSS.n8011 13.653
R10377 VSS.n8026 VSS.n8025 13.653
R10378 VSS.n8040 VSS.n8039 13.653
R10379 VSS.n8054 VSS.n8053 13.653
R10380 VSS.n8068 VSS.n8067 13.653
R10381 VSS.n8082 VSS.n8081 13.653
R10382 VSS.n8086 VSS.n8085 13.653
R10383 VSS.n8104 VSS.n8103 13.653
R10384 VSS.n8118 VSS.n8117 13.653
R10385 VSS.n8132 VSS.n8131 13.653
R10386 VSS.n8146 VSS.n8145 13.653
R10387 VSS.n8160 VSS.n8159 13.653
R10388 VSS.n8744 VSS.n8743 13.653
R10389 VSS.n8758 VSS.n8757 13.653
R10390 VSS.n8772 VSS.n8771 13.653
R10391 VSS.n8786 VSS.n8785 13.653
R10392 VSS.n8800 VSS.n8799 13.653
R10393 VSS.n8814 VSS.n8813 13.653
R10394 VSS.n8818 VSS.n8817 13.653
R10395 VSS.n8836 VSS.n8835 13.653
R10396 VSS.n8850 VSS.n8849 13.653
R10397 VSS.n8864 VSS.n8863 13.653
R10398 VSS.n8878 VSS.n8877 13.653
R10399 VSS.n8892 VSS.n8891 13.653
R10400 VSS.n8500 VSS.n8499 13.653
R10401 VSS.n8514 VSS.n8513 13.653
R10402 VSS.n8528 VSS.n8527 13.653
R10403 VSS.n8542 VSS.n8541 13.653
R10404 VSS.n8556 VSS.n8555 13.653
R10405 VSS.n8570 VSS.n8569 13.653
R10406 VSS.n8574 VSS.n8573 13.653
R10407 VSS.n8592 VSS.n8591 13.653
R10408 VSS.n8606 VSS.n8605 13.653
R10409 VSS.n8620 VSS.n8619 13.653
R10410 VSS.n8634 VSS.n8633 13.653
R10411 VSS.n8648 VSS.n8647 13.653
R10412 VSS.n9000 VSS.n8999 13.653
R10413 VSS.n9014 VSS.n9013 13.653
R10414 VSS.n9028 VSS.n9027 13.653
R10415 VSS.n9042 VSS.n9041 13.653
R10416 VSS.n9056 VSS.n9055 13.653
R10417 VSS.n9070 VSS.n9069 13.653
R10418 VSS.n9074 VSS.n9073 13.653
R10419 VSS.n9092 VSS.n9091 13.653
R10420 VSS.n9106 VSS.n9105 13.653
R10421 VSS.n9120 VSS.n9119 13.653
R10422 VSS.n9134 VSS.n9133 13.653
R10423 VSS.n9193 VSS.n9192 13.653
R10424 VSS.n5136 VSS.n1584 13.653
R10425 VSS.n5148 VSS.n1579 13.653
R10426 VSS.n5152 VSS.n1571 13.653
R10427 VSS.n5163 VSS.n1569 13.653
R10428 VSS.n5171 VSS.n1563 13.653
R10429 VSS.n5183 VSS.n1558 13.653
R10430 VSS.n5187 VSS.n1550 13.653
R10431 VSS.n5198 VSS.n1548 13.653
R10432 VSS.n5206 VSS.n1542 13.653
R10433 VSS.n5218 VSS.n1537 13.653
R10434 VSS.n5223 VSS.n1535 13.653
R10435 VSS.n5232 VSS.n1526 13.653
R10436 VSS.n5495 VSS.n1443 13.653
R10437 VSS.n5507 VSS.n1438 13.653
R10438 VSS.n5511 VSS.n1430 13.653
R10439 VSS.n5522 VSS.n1428 13.653
R10440 VSS.n5530 VSS.n1422 13.653
R10441 VSS.n5542 VSS.n1417 13.653
R10442 VSS.n5546 VSS.n1409 13.653
R10443 VSS.n5557 VSS.n1407 13.653
R10444 VSS.n5565 VSS.n1401 13.653
R10445 VSS.n5577 VSS.n1396 13.653
R10446 VSS.n5582 VSS.n1394 13.653
R10447 VSS.n5591 VSS.n1385 13.653
R10448 VSS.n5399 VSS.n5398 13.653
R10449 VSS.n5390 VSS.n5240 13.653
R10450 VSS.n5249 VSS.n5243 13.653
R10451 VSS.n5375 VSS.n5250 13.653
R10452 VSS.n5367 VSS.n5260 13.653
R10453 VSS.n5268 VSS.n5262 13.653
R10454 VSS.n5352 VSS.n5269 13.653
R10455 VSS.n5344 VSS.n5279 13.653
R10456 VSS.n5287 VSS.n5281 13.653
R10457 VSS.n5329 VSS.n5288 13.653
R10458 VSS.n5321 VSS.n5298 13.653
R10459 VSS.n5307 VSS.n5300 13.653
R10460 VSS.n781 VSS.n780 13.653
R10461 VSS.n793 VSS.n775 13.653
R10462 VSS.n797 VSS.n767 13.653
R10463 VSS.n808 VSS.n765 13.653
R10464 VSS.n816 VSS.n759 13.653
R10465 VSS.n828 VSS.n754 13.653
R10466 VSS.n832 VSS.n746 13.653
R10467 VSS.n843 VSS.n744 13.653
R10468 VSS.n851 VSS.n738 13.653
R10469 VSS.n863 VSS.n733 13.653
R10470 VSS.n867 VSS.n724 13.653
R10471 VSS.n878 VSS.n722 13.653
R10472 VSS.n5607 VSS.n5606 13.653
R10473 VSS.n5598 VSS.n523 13.653
R10474 VSS.n5777 VSS.n524 13.653
R10475 VSS.n5769 VSS.n534 13.653
R10476 VSS.n542 VSS.n536 13.653
R10477 VSS.n5754 VSS.n543 13.653
R10478 VSS.n5746 VSS.n553 13.653
R10479 VSS.n561 VSS.n555 13.653
R10480 VSS.n5731 VSS.n562 13.653
R10481 VSS.n5723 VSS.n572 13.653
R10482 VSS.n580 VSS.n574 13.653
R10483 VSS.n5708 VSS.n581 13.653
R10484 VSS.n920 VSS.n714 13.653
R10485 VSS.n928 VSS.n708 13.653
R10486 VSS.n940 VSS.n703 13.653
R10487 VSS.n944 VSS.n695 13.653
R10488 VSS.n955 VSS.n693 13.653
R10489 VSS.n963 VSS.n687 13.653
R10490 VSS.n975 VSS.n682 13.653
R10491 VSS.n979 VSS.n674 13.653
R10492 VSS.n990 VSS.n672 13.653
R10493 VSS.n998 VSS.n666 13.653
R10494 VSS.n1010 VSS.n661 13.653
R10495 VSS.n1014 VSS.n654 13.653
R10496 VSS.n1023 VSS.n1022 13.653
R10497 VSS.n1254 VSS.n1024 13.653
R10498 VSS.n1246 VSS.n1034 13.653
R10499 VSS.n1042 VSS.n1036 13.653
R10500 VSS.n1231 VSS.n1043 13.653
R10501 VSS.n1223 VSS.n1053 13.653
R10502 VSS.n1061 VSS.n1055 13.653
R10503 VSS.n1208 VSS.n1062 13.653
R10504 VSS.n1200 VSS.n1072 13.653
R10505 VSS.n1080 VSS.n1074 13.653
R10506 VSS.n1185 VSS.n1081 13.653
R10507 VSS.n1177 VSS.n1091 13.653
R10508 VSS.n3809 VSS.n3450 13.653
R10509 VSS.n3801 VSS.n3454 13.653
R10510 VSS.n3793 VSS.n3464 13.653
R10511 VSS.n3472 VSS.n3466 13.653
R10512 VSS.n3778 VSS.n3473 13.653
R10513 VSS.n3770 VSS.n3483 13.653
R10514 VSS.n3491 VSS.n3485 13.653
R10515 VSS.n3755 VSS.n3492 13.653
R10516 VSS.n3747 VSS.n3502 13.653
R10517 VSS.n3510 VSS.n3504 13.653
R10518 VSS.n3732 VSS.n3511 13.653
R10519 VSS.n3724 VSS.n3521 13.653
R10520 VSS.n3962 VSS.n3384 13.653
R10521 VSS.n3970 VSS.n3378 13.653
R10522 VSS.n3982 VSS.n3373 13.653
R10523 VSS.n3986 VSS.n3365 13.653
R10524 VSS.n3997 VSS.n3363 13.653
R10525 VSS.n4005 VSS.n3357 13.653
R10526 VSS.n4017 VSS.n3352 13.653
R10527 VSS.n4021 VSS.n3344 13.653
R10528 VSS.n4032 VSS.n3342 13.653
R10529 VSS.n4040 VSS.n3336 13.653
R10530 VSS.n4052 VSS.n3331 13.653
R10531 VSS.n4056 VSS.n3324 13.653
R10532 VSS.n3565 VSS.n3562 13.653
R10533 VSS.n3708 VSS.n3563 13.653
R10534 VSS.n3700 VSS.n3576 13.653
R10535 VSS.n3584 VSS.n3578 13.653
R10536 VSS.n3685 VSS.n3585 13.653
R10537 VSS.n3677 VSS.n3595 13.653
R10538 VSS.n3603 VSS.n3597 13.653
R10539 VSS.n3662 VSS.n3604 13.653
R10540 VSS.n3654 VSS.n3614 13.653
R10541 VSS.n3622 VSS.n3616 13.653
R10542 VSS.n3639 VSS.n3623 13.653
R10543 VSS.n3629 VSS.n3387 13.653
R10544 VSS.n4177 VSS.n4174 13.653
R10545 VSS.n4312 VSS.n4175 13.653
R10546 VSS.n4304 VSS.n4188 13.653
R10547 VSS.n4196 VSS.n4190 13.653
R10548 VSS.n4289 VSS.n4197 13.653
R10549 VSS.n4281 VSS.n4207 13.653
R10550 VSS.n4215 VSS.n4209 13.653
R10551 VSS.n4266 VSS.n4216 13.653
R10552 VSS.n4258 VSS.n4226 13.653
R10553 VSS.n4234 VSS.n4228 13.653
R10554 VSS.n4243 VSS.n4235 13.653
R10555 VSS.n4535 VSS.n3226 13.653
R10556 VSS.n4065 VSS.n4064 13.653
R10557 VSS.n4405 VSS.n4066 13.653
R10558 VSS.n4397 VSS.n4076 13.653
R10559 VSS.n4084 VSS.n4078 13.653
R10560 VSS.n4382 VSS.n4085 13.653
R10561 VSS.n4374 VSS.n4095 13.653
R10562 VSS.n4103 VSS.n4097 13.653
R10563 VSS.n4359 VSS.n4104 13.653
R10564 VSS.n4351 VSS.n4114 13.653
R10565 VSS.n4122 VSS.n4116 13.653
R10566 VSS.n4336 VSS.n4123 13.653
R10567 VSS.n4328 VSS.n4133 13.653
R10568 VSS.n4655 VSS.n4653 13.653
R10569 VSS.n5014 VSS.n4654 13.653
R10570 VSS.n5006 VSS.n4666 13.653
R10571 VSS.n4674 VSS.n4668 13.653
R10572 VSS.n4991 VSS.n4675 13.653
R10573 VSS.n4983 VSS.n4685 13.653
R10574 VSS.n4693 VSS.n4687 13.653
R10575 VSS.n4968 VSS.n4694 13.653
R10576 VSS.n4960 VSS.n4704 13.653
R10577 VSS.n4712 VSS.n4706 13.653
R10578 VSS.n4945 VSS.n4713 13.653
R10579 VSS.n4937 VSS.n4723 13.653
R10580 VSS.n4548 VSS.n3217 13.653
R10581 VSS.n4552 VSS.n3209 13.653
R10582 VSS.n4563 VSS.n3207 13.653
R10583 VSS.n4571 VSS.n3201 13.653
R10584 VSS.n4583 VSS.n3196 13.653
R10585 VSS.n4587 VSS.n3188 13.653
R10586 VSS.n4598 VSS.n3186 13.653
R10587 VSS.n4606 VSS.n3180 13.653
R10588 VSS.n4618 VSS.n3175 13.653
R10589 VSS.n4622 VSS.n3167 13.653
R10590 VSS.n4633 VSS.n3165 13.653
R10591 VSS.n4641 VSS.n3159 13.653
R10592 VSS.n4767 VSS.n4764 13.653
R10593 VSS.n4921 VSS.n4765 13.653
R10594 VSS.n4913 VSS.n4778 13.653
R10595 VSS.n4786 VSS.n4780 13.653
R10596 VSS.n4898 VSS.n4787 13.653
R10597 VSS.n4890 VSS.n4797 13.653
R10598 VSS.n4805 VSS.n4799 13.653
R10599 VSS.n4875 VSS.n4806 13.653
R10600 VSS.n4867 VSS.n4816 13.653
R10601 VSS.n4824 VSS.n4818 13.653
R10602 VSS.n4852 VSS.n4825 13.653
R10603 VSS.n4844 VSS.n4835 13.653
R10604 VSS.n384 VSS.n383 13.552
R10605 VSS.n391 VSS.n390 13.552
R10606 VSS.n393 VSS.n363 13.552
R10607 VSS.n415 VSS.n414 13.552
R10608 VSS.n422 VSS.n421 13.552
R10609 VSS.n430 VSS.n429 13.552
R10610 VSS.n18176 VSS.n18175 13.552
R10611 VSS.n18183 VSS.n18182 13.552
R10612 VSS.n18185 VSS.n18155 13.552
R10613 VSS.n18207 VSS.n18206 13.552
R10614 VSS.n18145 VSS.n18142 13.552
R10615 VSS.n18221 VSS.n18220 13.552
R10616 VSS.n17949 VSS.n17948 13.511
R10617 VSS.n10579 VSS 13.314
R10618 VSS.n17856 VSS.n17805 13.058
R10619 VSS.n17436 VSS.n17435 13.014
R10620 VSS.n17268 VSS.n17267 13.014
R10621 VSS.n17100 VSS.n17099 13.014
R10622 VSS.n16932 VSS.n16931 13.014
R10623 VSS.n16764 VSS.n16763 13.014
R10624 VSS.n16596 VSS.n16595 13.014
R10625 VSS.n10401 VSS.n10400 13.014
R10626 VSS.n6247 VSS.n6107 13.014
R10627 VSS.n6311 VSS.n5991 13.014
R10628 VSS.n6375 VSS.n5875 13.014
R10629 VSS.n5837 VSS.n5831 13.014
R10630 VSS VSS.n17984 12.977
R10631 VSS.n386 VSS.n367 12.413
R10632 VSS.n426 VSS.n349 12.413
R10633 VSS.n18178 VSS.n18159 12.413
R10634 VSS.n18214 VSS.n18139 12.413
R10635 VSS.n17880 VSS.n17793 12.412
R10636 VSS.n14317 VSS.n14316 11.666
R10637 VSS.n14329 VSS.n14328 11.666
R10638 VSS.n14341 VSS.n14340 11.666
R10639 VSS.n14353 VSS.n14352 11.666
R10640 VSS.n14365 VSS.n14364 11.666
R10641 VSS.n14377 VSS.n14376 11.666
R10642 VSS.n14389 VSS.n14388 11.666
R10643 VSS.n14401 VSS.n14400 11.666
R10644 VSS.n14413 VSS.n14412 11.666
R10645 VSS.n14137 VSS.n14136 11.666
R10646 VSS.n14149 VSS.n14148 11.666
R10647 VSS.n14161 VSS.n14160 11.666
R10648 VSS.n14173 VSS.n14172 11.666
R10649 VSS.n14185 VSS.n14184 11.666
R10650 VSS.n14197 VSS.n14196 11.666
R10651 VSS.n14209 VSS.n14208 11.666
R10652 VSS.n14221 VSS.n14220 11.666
R10653 VSS.n14233 VSS.n14232 11.666
R10654 VSS.n17519 VSS.n17518 11.666
R10655 VSS.n17507 VSS.n17506 11.666
R10656 VSS.n17495 VSS.n17494 11.666
R10657 VSS.n17483 VSS.n17482 11.666
R10658 VSS.n17474 VSS.n17473 11.666
R10659 VSS.n17459 VSS.n17458 11.666
R10660 VSS.n17447 VSS.n17446 11.666
R10661 VSS.n17435 VSS.n17434 11.666
R10662 VSS.n17351 VSS.n17350 11.666
R10663 VSS.n17339 VSS.n17338 11.666
R10664 VSS.n17327 VSS.n17326 11.666
R10665 VSS.n17315 VSS.n17314 11.666
R10666 VSS.n17306 VSS.n17305 11.666
R10667 VSS.n17291 VSS.n17290 11.666
R10668 VSS.n17279 VSS.n17278 11.666
R10669 VSS.n17267 VSS.n17266 11.666
R10670 VSS.n17183 VSS.n17182 11.666
R10671 VSS.n17171 VSS.n17170 11.666
R10672 VSS.n17159 VSS.n17158 11.666
R10673 VSS.n17147 VSS.n17146 11.666
R10674 VSS.n17138 VSS.n17137 11.666
R10675 VSS.n17123 VSS.n17122 11.666
R10676 VSS.n17111 VSS.n17110 11.666
R10677 VSS.n17099 VSS.n17098 11.666
R10678 VSS.n17015 VSS.n17014 11.666
R10679 VSS.n17003 VSS.n17002 11.666
R10680 VSS.n16991 VSS.n16990 11.666
R10681 VSS.n16979 VSS.n16978 11.666
R10682 VSS.n16970 VSS.n16969 11.666
R10683 VSS.n16955 VSS.n16954 11.666
R10684 VSS.n16943 VSS.n16942 11.666
R10685 VSS.n16931 VSS.n16930 11.666
R10686 VSS.n16847 VSS.n16846 11.666
R10687 VSS.n16835 VSS.n16834 11.666
R10688 VSS.n16823 VSS.n16822 11.666
R10689 VSS.n16811 VSS.n16810 11.666
R10690 VSS.n16802 VSS.n16801 11.666
R10691 VSS.n16787 VSS.n16786 11.666
R10692 VSS.n16775 VSS.n16774 11.666
R10693 VSS.n16763 VSS.n16762 11.666
R10694 VSS.n16679 VSS.n16678 11.666
R10695 VSS.n16667 VSS.n16666 11.666
R10696 VSS.n16655 VSS.n16654 11.666
R10697 VSS.n16643 VSS.n16642 11.666
R10698 VSS.n16634 VSS.n16633 11.666
R10699 VSS.n16619 VSS.n16618 11.666
R10700 VSS.n16607 VSS.n16606 11.666
R10701 VSS.n16595 VSS.n16594 11.666
R10702 VSS.n13914 VSS.n13913 11.666
R10703 VSS.n13926 VSS.n13925 11.666
R10704 VSS.n13938 VSS.n13937 11.666
R10705 VSS.n13950 VSS.n13949 11.666
R10706 VSS.n13962 VSS.n13961 11.666
R10707 VSS.n13974 VSS.n13973 11.666
R10708 VSS.n13986 VSS.n13985 11.666
R10709 VSS.n13998 VSS.n13997 11.666
R10710 VSS.n14010 VSS.n14009 11.666
R10711 VSS.n13734 VSS.n13733 11.666
R10712 VSS.n13746 VSS.n13745 11.666
R10713 VSS.n13758 VSS.n13757 11.666
R10714 VSS.n13770 VSS.n13769 11.666
R10715 VSS.n13782 VSS.n13781 11.666
R10716 VSS.n13794 VSS.n13793 11.666
R10717 VSS.n13806 VSS.n13805 11.666
R10718 VSS.n13818 VSS.n13817 11.666
R10719 VSS.n13830 VSS.n13829 11.666
R10720 VSS.n13554 VSS.n13553 11.666
R10721 VSS.n13566 VSS.n13565 11.666
R10722 VSS.n13578 VSS.n13577 11.666
R10723 VSS.n13590 VSS.n13589 11.666
R10724 VSS.n13602 VSS.n13601 11.666
R10725 VSS.n13614 VSS.n13613 11.666
R10726 VSS.n13626 VSS.n13625 11.666
R10727 VSS.n13638 VSS.n13637 11.666
R10728 VSS.n13650 VSS.n13649 11.666
R10729 VSS.n13374 VSS.n13373 11.666
R10730 VSS.n13386 VSS.n13385 11.666
R10731 VSS.n13398 VSS.n13397 11.666
R10732 VSS.n13410 VSS.n13409 11.666
R10733 VSS.n13422 VSS.n13421 11.666
R10734 VSS.n13434 VSS.n13433 11.666
R10735 VSS.n13446 VSS.n13445 11.666
R10736 VSS.n13458 VSS.n13457 11.666
R10737 VSS.n13470 VSS.n13469 11.666
R10738 VSS.n13194 VSS.n13193 11.666
R10739 VSS.n13206 VSS.n13205 11.666
R10740 VSS.n13218 VSS.n13217 11.666
R10741 VSS.n13230 VSS.n13229 11.666
R10742 VSS.n13242 VSS.n13241 11.666
R10743 VSS.n13254 VSS.n13253 11.666
R10744 VSS.n13266 VSS.n13265 11.666
R10745 VSS.n13278 VSS.n13277 11.666
R10746 VSS.n13290 VSS.n13289 11.666
R10747 VSS.n13014 VSS.n13013 11.666
R10748 VSS.n13026 VSS.n13025 11.666
R10749 VSS.n13038 VSS.n13037 11.666
R10750 VSS.n13050 VSS.n13049 11.666
R10751 VSS.n13062 VSS.n13061 11.666
R10752 VSS.n13074 VSS.n13073 11.666
R10753 VSS.n13086 VSS.n13085 11.666
R10754 VSS.n13098 VSS.n13097 11.666
R10755 VSS.n13110 VSS.n13109 11.666
R10756 VSS.n12834 VSS.n12833 11.666
R10757 VSS.n12846 VSS.n12845 11.666
R10758 VSS.n12858 VSS.n12857 11.666
R10759 VSS.n12870 VSS.n12869 11.666
R10760 VSS.n12882 VSS.n12881 11.666
R10761 VSS.n12894 VSS.n12893 11.666
R10762 VSS.n12906 VSS.n12905 11.666
R10763 VSS.n12918 VSS.n12917 11.666
R10764 VSS.n12930 VSS.n12929 11.666
R10765 VSS.n12654 VSS.n12653 11.666
R10766 VSS.n12666 VSS.n12665 11.666
R10767 VSS.n12678 VSS.n12677 11.666
R10768 VSS.n12690 VSS.n12689 11.666
R10769 VSS.n12702 VSS.n12701 11.666
R10770 VSS.n12714 VSS.n12713 11.666
R10771 VSS.n12726 VSS.n12725 11.666
R10772 VSS.n12738 VSS.n12737 11.666
R10773 VSS.n12750 VSS.n12749 11.666
R10774 VSS.n9321 VSS.n9320 11.666
R10775 VSS.n9309 VSS.n9308 11.666
R10776 VSS.n9297 VSS.n9296 11.666
R10777 VSS.n9285 VSS.n9284 11.666
R10778 VSS.n9273 VSS.n9272 11.666
R10779 VSS.n9264 VSS.n9263 11.666
R10780 VSS.n9249 VSS.n9248 11.666
R10781 VSS.n9237 VSS.n9236 11.666
R10782 VSS.n9225 VSS.n9224 11.666
R10783 VSS.n9489 VSS.n9488 11.666
R10784 VSS.n9477 VSS.n9476 11.666
R10785 VSS.n9465 VSS.n9464 11.666
R10786 VSS.n9453 VSS.n9452 11.666
R10787 VSS.n9441 VSS.n9440 11.666
R10788 VSS.n9432 VSS.n9431 11.666
R10789 VSS.n9417 VSS.n9416 11.666
R10790 VSS.n9405 VSS.n9404 11.666
R10791 VSS.n9393 VSS.n9392 11.666
R10792 VSS.n9657 VSS.n9656 11.666
R10793 VSS.n9645 VSS.n9644 11.666
R10794 VSS.n9633 VSS.n9632 11.666
R10795 VSS.n9621 VSS.n9620 11.666
R10796 VSS.n9609 VSS.n9608 11.666
R10797 VSS.n9600 VSS.n9599 11.666
R10798 VSS.n9585 VSS.n9584 11.666
R10799 VSS.n9573 VSS.n9572 11.666
R10800 VSS.n9561 VSS.n9560 11.666
R10801 VSS.n9825 VSS.n9824 11.666
R10802 VSS.n9813 VSS.n9812 11.666
R10803 VSS.n9801 VSS.n9800 11.666
R10804 VSS.n9789 VSS.n9788 11.666
R10805 VSS.n9777 VSS.n9776 11.666
R10806 VSS.n9768 VSS.n9767 11.666
R10807 VSS.n9753 VSS.n9752 11.666
R10808 VSS.n9741 VSS.n9740 11.666
R10809 VSS.n9729 VSS.n9728 11.666
R10810 VSS.n9993 VSS.n9992 11.666
R10811 VSS.n9981 VSS.n9980 11.666
R10812 VSS.n9969 VSS.n9968 11.666
R10813 VSS.n9957 VSS.n9956 11.666
R10814 VSS.n9945 VSS.n9944 11.666
R10815 VSS.n9936 VSS.n9935 11.666
R10816 VSS.n9921 VSS.n9920 11.666
R10817 VSS.n9909 VSS.n9908 11.666
R10818 VSS.n9897 VSS.n9896 11.666
R10819 VSS.n10161 VSS.n10160 11.666
R10820 VSS.n10149 VSS.n10148 11.666
R10821 VSS.n10137 VSS.n10136 11.666
R10822 VSS.n10125 VSS.n10124 11.666
R10823 VSS.n10113 VSS.n10112 11.666
R10824 VSS.n10104 VSS.n10103 11.666
R10825 VSS.n10089 VSS.n10088 11.666
R10826 VSS.n10077 VSS.n10076 11.666
R10827 VSS.n10065 VSS.n10064 11.666
R10828 VSS.n10329 VSS.n10328 11.666
R10829 VSS.n10317 VSS.n10316 11.666
R10830 VSS.n10305 VSS.n10304 11.666
R10831 VSS.n10293 VSS.n10292 11.666
R10832 VSS.n10281 VSS.n10280 11.666
R10833 VSS.n10272 VSS.n10271 11.666
R10834 VSS.n10257 VSS.n10256 11.666
R10835 VSS.n10245 VSS.n10244 11.666
R10836 VSS.n10233 VSS.n10232 11.666
R10837 VSS.n10484 VSS.n10483 11.666
R10838 VSS.n10472 VSS.n10471 11.666
R10839 VSS.n10460 VSS.n10459 11.666
R10840 VSS.n10448 VSS.n10447 11.666
R10841 VSS.n10439 VSS.n10438 11.666
R10842 VSS.n10424 VSS.n10423 11.666
R10843 VSS.n10412 VSS.n10411 11.666
R10844 VSS.n10400 VSS.n10399 11.666
R10845 VSS.n2456 VSS.n2306 11.666
R10846 VSS.n2446 VSS.n2310 11.666
R10847 VSS.n2386 VSS.n2305 11.666
R10848 VSS.n2389 VSS.n2311 11.666
R10849 VSS.n2393 VSS.n2304 11.666
R10850 VSS.n2459 VSS.n2312 11.666
R10851 VSS.n2399 VSS.n2308 11.666
R10852 VSS.n2406 VSS.n2405 11.666
R10853 VSS.n2546 VSS.n2216 11.666
R10854 VSS.n2536 VSS.n2220 11.666
R10855 VSS.n2476 VSS.n2215 11.666
R10856 VSS.n2479 VSS.n2221 11.666
R10857 VSS.n2483 VSS.n2214 11.666
R10858 VSS.n2549 VSS.n2222 11.666
R10859 VSS.n2489 VSS.n2218 11.666
R10860 VSS.n2496 VSS.n2495 11.666
R10861 VSS.n2636 VSS.n2126 11.666
R10862 VSS.n2626 VSS.n2130 11.666
R10863 VSS.n2566 VSS.n2125 11.666
R10864 VSS.n2569 VSS.n2131 11.666
R10865 VSS.n2573 VSS.n2124 11.666
R10866 VSS.n2639 VSS.n2132 11.666
R10867 VSS.n2579 VSS.n2128 11.666
R10868 VSS.n2586 VSS.n2585 11.666
R10869 VSS.n2726 VSS.n2036 11.666
R10870 VSS.n2716 VSS.n2040 11.666
R10871 VSS.n2656 VSS.n2035 11.666
R10872 VSS.n2659 VSS.n2041 11.666
R10873 VSS.n2663 VSS.n2034 11.666
R10874 VSS.n2729 VSS.n2042 11.666
R10875 VSS.n2669 VSS.n2038 11.666
R10876 VSS.n2676 VSS.n2675 11.666
R10877 VSS.n2816 VSS.n1946 11.666
R10878 VSS.n2806 VSS.n1950 11.666
R10879 VSS.n2746 VSS.n1945 11.666
R10880 VSS.n2749 VSS.n1951 11.666
R10881 VSS.n2753 VSS.n1944 11.666
R10882 VSS.n2819 VSS.n1952 11.666
R10883 VSS.n2759 VSS.n1948 11.666
R10884 VSS.n2766 VSS.n2765 11.666
R10885 VSS.n2906 VSS.n1856 11.666
R10886 VSS.n2896 VSS.n1860 11.666
R10887 VSS.n2836 VSS.n1855 11.666
R10888 VSS.n2839 VSS.n1861 11.666
R10889 VSS.n2843 VSS.n1854 11.666
R10890 VSS.n2909 VSS.n1862 11.666
R10891 VSS.n2849 VSS.n1858 11.666
R10892 VSS.n2856 VSS.n2855 11.666
R10893 VSS.n2996 VSS.n1766 11.666
R10894 VSS.n2986 VSS.n1770 11.666
R10895 VSS.n2926 VSS.n1765 11.666
R10896 VSS.n2929 VSS.n1771 11.666
R10897 VSS.n2933 VSS.n1764 11.666
R10898 VSS.n2999 VSS.n1772 11.666
R10899 VSS.n2939 VSS.n1768 11.666
R10900 VSS.n2946 VSS.n2945 11.666
R10901 VSS.n3086 VSS.n1676 11.666
R10902 VSS.n3076 VSS.n1680 11.666
R10903 VSS.n3016 VSS.n1675 11.666
R10904 VSS.n3019 VSS.n1681 11.666
R10905 VSS.n3023 VSS.n1674 11.666
R10906 VSS.n3089 VSS.n1682 11.666
R10907 VSS.n3029 VSS.n1678 11.666
R10908 VSS.n3036 VSS.n3035 11.666
R10909 VSS.n6129 VSS.n6081 11.666
R10910 VSS.n6137 VSS.n6080 11.666
R10911 VSS.n6145 VSS.n6082 11.666
R10912 VSS.n6153 VSS.n6079 11.666
R10913 VSS.n6161 VSS.n6083 11.666
R10914 VSS.n6169 VSS.n6078 11.666
R10915 VSS.n6177 VSS.n6084 11.666
R10916 VSS.n6185 VSS.n6107 11.666
R10917 VSS.n6013 VSS.n5965 11.666
R10918 VSS.n6021 VSS.n5964 11.666
R10919 VSS.n6029 VSS.n5966 11.666
R10920 VSS.n6037 VSS.n5963 11.666
R10921 VSS.n6045 VSS.n5967 11.666
R10922 VSS.n6053 VSS.n5962 11.666
R10923 VSS.n6061 VSS.n5968 11.666
R10924 VSS.n6069 VSS.n5991 11.666
R10925 VSS.n5897 VSS.n5849 11.666
R10926 VSS.n5905 VSS.n5848 11.666
R10927 VSS.n5913 VSS.n5850 11.666
R10928 VSS.n5921 VSS.n5847 11.666
R10929 VSS.n5929 VSS.n5851 11.666
R10930 VSS.n5937 VSS.n5846 11.666
R10931 VSS.n5945 VSS.n5852 11.666
R10932 VSS.n5953 VSS.n5875 11.666
R10933 VSS.n7040 VSS.n5790 11.666
R10934 VSS.n7034 VSS.n5795 11.666
R10935 VSS.n7028 VSS.n5801 11.666
R10936 VSS.n7022 VSS.n5807 11.666
R10937 VSS.n7016 VSS.n5813 11.666
R10938 VSS.n7010 VSS.n5818 11.666
R10939 VSS.n7004 VSS.n5825 11.666
R10940 VSS.n6998 VSS.n5831 11.666
R10941 VSS.n6851 VSS.n6429 11.666
R10942 VSS.n6929 VSS.n6423 11.666
R10943 VSS.n6919 VSS.n6420 11.666
R10944 VSS.n6860 VSS.n6424 11.666
R10945 VSS.n6863 VSS.n6419 11.666
R10946 VSS.n6867 VSS.n6425 11.666
R10947 VSS.n6871 VSS.n6418 11.666
R10948 VSS.n6933 VSS.n6426 11.666
R10949 VSS.n6877 VSS.n6422 11.666
R10950 VSS.n6761 VSS.n6519 11.666
R10951 VSS.n6839 VSS.n6513 11.666
R10952 VSS.n6829 VSS.n6510 11.666
R10953 VSS.n6770 VSS.n6514 11.666
R10954 VSS.n6773 VSS.n6509 11.666
R10955 VSS.n6777 VSS.n6515 11.666
R10956 VSS.n6781 VSS.n6508 11.666
R10957 VSS.n6843 VSS.n6516 11.666
R10958 VSS.n6787 VSS.n6512 11.666
R10959 VSS.n6671 VSS.n6609 11.666
R10960 VSS.n6749 VSS.n6603 11.666
R10961 VSS.n6739 VSS.n6600 11.666
R10962 VSS.n6680 VSS.n6604 11.666
R10963 VSS.n6683 VSS.n6599 11.666
R10964 VSS.n6687 VSS.n6605 11.666
R10965 VSS.n6691 VSS.n6598 11.666
R10966 VSS.n6753 VSS.n6606 11.666
R10967 VSS.n6697 VSS.n6602 11.666
R10968 VSS.n14641 VSS.n14638 11.636
R10969 VSS.n14638 VSS.n14635 11.636
R10970 VSS.n14635 VSS.n14632 11.636
R10971 VSS.n14632 VSS.n14629 11.636
R10972 VSS.n14629 VSS.n14626 11.636
R10973 VSS.n14626 VSS.n14623 11.636
R10974 VSS.n14623 VSS.n14620 11.636
R10975 VSS.n14620 VSS.n14617 11.636
R10976 VSS.n14617 VSS.n14614 11.636
R10977 VSS.n14614 VSS.n14611 11.636
R10978 VSS.n14611 VSS.n14608 11.636
R10979 VSS.n16569 VSS.n16566 11.636
R10980 VSS.n16566 VSS.n16563 11.636
R10981 VSS.n16563 VSS.n16560 11.636
R10982 VSS.n16560 VSS.n16557 11.636
R10983 VSS.n16557 VSS.n16554 11.636
R10984 VSS.n16554 VSS.n16551 11.636
R10985 VSS.n16551 VSS.n16548 11.636
R10986 VSS.n16548 VSS.n16545 11.636
R10987 VSS.n16545 VSS.n16542 11.636
R10988 VSS.n16542 VSS.n16539 11.636
R10989 VSS.n16539 VSS.n16536 11.636
R10990 VSS.n16317 VSS.n16314 11.636
R10991 VSS.n16314 VSS.n16311 11.636
R10992 VSS.n16311 VSS.n16308 11.636
R10993 VSS.n16308 VSS.n16305 11.636
R10994 VSS.n16305 VSS.n16302 11.636
R10995 VSS.n16302 VSS.n16299 11.636
R10996 VSS.n16299 VSS.n16296 11.636
R10997 VSS.n16296 VSS.n16293 11.636
R10998 VSS.n16293 VSS.n16290 11.636
R10999 VSS.n16533 VSS.n16530 11.636
R11000 VSS.n16062 VSS.n16059 11.636
R11001 VSS.n16059 VSS.n16056 11.636
R11002 VSS.n16056 VSS.n16053 11.636
R11003 VSS.n16053 VSS.n16050 11.636
R11004 VSS.n16050 VSS.n16047 11.636
R11005 VSS.n16323 VSS.n16320 11.636
R11006 VSS.n16326 VSS.n16323 11.636
R11007 VSS.n16329 VSS.n16326 11.636
R11008 VSS.n16332 VSS.n16329 11.636
R11009 VSS.n16333 VSS.n16332 11.636
R11010 VSS.n15817 VSS.n15814 11.636
R11011 VSS.n15814 VSS.n15811 11.636
R11012 VSS.n15811 VSS.n15808 11.636
R11013 VSS.n15808 VSS.n15805 11.636
R11014 VSS.n15805 VSS.n15802 11.636
R11015 VSS.n16068 VSS.n16065 11.636
R11016 VSS.n16071 VSS.n16068 11.636
R11017 VSS.n16074 VSS.n16071 11.636
R11018 VSS.n16077 VSS.n16074 11.636
R11019 VSS.n16078 VSS.n16077 11.636
R11020 VSS.n15574 VSS.n15571 11.636
R11021 VSS.n15571 VSS.n15568 11.636
R11022 VSS.n15568 VSS.n15565 11.636
R11023 VSS.n15565 VSS.n15562 11.636
R11024 VSS.n15562 VSS.n15559 11.636
R11025 VSS.n15823 VSS.n15820 11.636
R11026 VSS.n15826 VSS.n15823 11.636
R11027 VSS.n15829 VSS.n15826 11.636
R11028 VSS.n15832 VSS.n15829 11.636
R11029 VSS.n15833 VSS.n15832 11.636
R11030 VSS.n15329 VSS.n15326 11.636
R11031 VSS.n15326 VSS.n15323 11.636
R11032 VSS.n15323 VSS.n15320 11.636
R11033 VSS.n15320 VSS.n15317 11.636
R11034 VSS.n15317 VSS.n15314 11.636
R11035 VSS.n15580 VSS.n15577 11.636
R11036 VSS.n15583 VSS.n15580 11.636
R11037 VSS.n15586 VSS.n15583 11.636
R11038 VSS.n15589 VSS.n15586 11.636
R11039 VSS.n15590 VSS.n15589 11.636
R11040 VSS.n15086 VSS.n15083 11.636
R11041 VSS.n15083 VSS.n15080 11.636
R11042 VSS.n15080 VSS.n15077 11.636
R11043 VSS.n15077 VSS.n15074 11.636
R11044 VSS.n15074 VSS.n15071 11.636
R11045 VSS.n15335 VSS.n15332 11.636
R11046 VSS.n15338 VSS.n15335 11.636
R11047 VSS.n15341 VSS.n15338 11.636
R11048 VSS.n15344 VSS.n15341 11.636
R11049 VSS.n15345 VSS.n15344 11.636
R11050 VSS.n14829 VSS.n14826 11.636
R11051 VSS.n14826 VSS.n14823 11.636
R11052 VSS.n14823 VSS.n14820 11.636
R11053 VSS.n14820 VSS.n14817 11.636
R11054 VSS.n14817 VSS.n14814 11.636
R11055 VSS.n15092 VSS.n15089 11.636
R11056 VSS.n15095 VSS.n15092 11.636
R11057 VSS.n15098 VSS.n15095 11.636
R11058 VSS.n15101 VSS.n15098 11.636
R11059 VSS.n15102 VSS.n15101 11.636
R11060 VSS.n14605 VSS.n14602 11.636
R11061 VSS.n14835 VSS.n14832 11.636
R11062 VSS.n14838 VSS.n14835 11.636
R11063 VSS.n14841 VSS.n14838 11.636
R11064 VSS.n14844 VSS.n14841 11.636
R11065 VSS.n14847 VSS.n14844 11.636
R11066 VSS.n14850 VSS.n14847 11.636
R11067 VSS.n14853 VSS.n14850 11.636
R11068 VSS.n14856 VSS.n14853 11.636
R11069 VSS.n14857 VSS.n14856 11.636
R11070 VSS.n10690 VSS.n10687 11.636
R11071 VSS.n10687 VSS.n10684 11.636
R11072 VSS.n10684 VSS.n10681 11.636
R11073 VSS.n10681 VSS.n10678 11.636
R11074 VSS.n10678 VSS.n10675 11.636
R11075 VSS.n10675 VSS.n10672 11.636
R11076 VSS.n10672 VSS.n10669 11.636
R11077 VSS.n10669 VSS.n10666 11.636
R11078 VSS.n10666 VSS.n10663 11.636
R11079 VSS.n10663 VSS.n10660 11.636
R11080 VSS.n10660 VSS.n10657 11.636
R11081 VSS.n12618 VSS.n12615 11.636
R11082 VSS.n12615 VSS.n12612 11.636
R11083 VSS.n12612 VSS.n12609 11.636
R11084 VSS.n12609 VSS.n12606 11.636
R11085 VSS.n12606 VSS.n12603 11.636
R11086 VSS.n12603 VSS.n12600 11.636
R11087 VSS.n12600 VSS.n12597 11.636
R11088 VSS.n12597 VSS.n12594 11.636
R11089 VSS.n12594 VSS.n12591 11.636
R11090 VSS.n12591 VSS.n12588 11.636
R11091 VSS.n12588 VSS.n12585 11.636
R11092 VSS.n12366 VSS.n12363 11.636
R11093 VSS.n12363 VSS.n12360 11.636
R11094 VSS.n12360 VSS.n12357 11.636
R11095 VSS.n12357 VSS.n12354 11.636
R11096 VSS.n12354 VSS.n12351 11.636
R11097 VSS.n12351 VSS.n12348 11.636
R11098 VSS.n12348 VSS.n12345 11.636
R11099 VSS.n12345 VSS.n12342 11.636
R11100 VSS.n12342 VSS.n12339 11.636
R11101 VSS.n12582 VSS.n12579 11.636
R11102 VSS.n12111 VSS.n12108 11.636
R11103 VSS.n12108 VSS.n12105 11.636
R11104 VSS.n12105 VSS.n12102 11.636
R11105 VSS.n12102 VSS.n12099 11.636
R11106 VSS.n12099 VSS.n12096 11.636
R11107 VSS.n12372 VSS.n12369 11.636
R11108 VSS.n12375 VSS.n12372 11.636
R11109 VSS.n12378 VSS.n12375 11.636
R11110 VSS.n12381 VSS.n12378 11.636
R11111 VSS.n12382 VSS.n12381 11.636
R11112 VSS.n11866 VSS.n11863 11.636
R11113 VSS.n11863 VSS.n11860 11.636
R11114 VSS.n11860 VSS.n11857 11.636
R11115 VSS.n11857 VSS.n11854 11.636
R11116 VSS.n11854 VSS.n11851 11.636
R11117 VSS.n12117 VSS.n12114 11.636
R11118 VSS.n12120 VSS.n12117 11.636
R11119 VSS.n12123 VSS.n12120 11.636
R11120 VSS.n12126 VSS.n12123 11.636
R11121 VSS.n12127 VSS.n12126 11.636
R11122 VSS.n11623 VSS.n11620 11.636
R11123 VSS.n11620 VSS.n11617 11.636
R11124 VSS.n11617 VSS.n11614 11.636
R11125 VSS.n11614 VSS.n11611 11.636
R11126 VSS.n11611 VSS.n11608 11.636
R11127 VSS.n11872 VSS.n11869 11.636
R11128 VSS.n11875 VSS.n11872 11.636
R11129 VSS.n11878 VSS.n11875 11.636
R11130 VSS.n11881 VSS.n11878 11.636
R11131 VSS.n11882 VSS.n11881 11.636
R11132 VSS.n11378 VSS.n11375 11.636
R11133 VSS.n11375 VSS.n11372 11.636
R11134 VSS.n11372 VSS.n11369 11.636
R11135 VSS.n11369 VSS.n11366 11.636
R11136 VSS.n11366 VSS.n11363 11.636
R11137 VSS.n11629 VSS.n11626 11.636
R11138 VSS.n11632 VSS.n11629 11.636
R11139 VSS.n11635 VSS.n11632 11.636
R11140 VSS.n11638 VSS.n11635 11.636
R11141 VSS.n11639 VSS.n11638 11.636
R11142 VSS.n11135 VSS.n11132 11.636
R11143 VSS.n11132 VSS.n11129 11.636
R11144 VSS.n11129 VSS.n11126 11.636
R11145 VSS.n11126 VSS.n11123 11.636
R11146 VSS.n11123 VSS.n11120 11.636
R11147 VSS.n11384 VSS.n11381 11.636
R11148 VSS.n11387 VSS.n11384 11.636
R11149 VSS.n11390 VSS.n11387 11.636
R11150 VSS.n11393 VSS.n11390 11.636
R11151 VSS.n11394 VSS.n11393 11.636
R11152 VSS.n10878 VSS.n10875 11.636
R11153 VSS.n10875 VSS.n10872 11.636
R11154 VSS.n10872 VSS.n10869 11.636
R11155 VSS.n10869 VSS.n10866 11.636
R11156 VSS.n10866 VSS.n10863 11.636
R11157 VSS.n11141 VSS.n11138 11.636
R11158 VSS.n11144 VSS.n11141 11.636
R11159 VSS.n11147 VSS.n11144 11.636
R11160 VSS.n11150 VSS.n11147 11.636
R11161 VSS.n11151 VSS.n11150 11.636
R11162 VSS.n10654 VSS.n10651 11.636
R11163 VSS.n10884 VSS.n10881 11.636
R11164 VSS.n10887 VSS.n10884 11.636
R11165 VSS.n10890 VSS.n10887 11.636
R11166 VSS.n10893 VSS.n10890 11.636
R11167 VSS.n10896 VSS.n10893 11.636
R11168 VSS.n10899 VSS.n10896 11.636
R11169 VSS.n10902 VSS.n10899 11.636
R11170 VSS.n10905 VSS.n10902 11.636
R11171 VSS.n10906 VSS.n10905 11.636
R11172 VSS.n7258 VSS.n7255 11.636
R11173 VSS.n7255 VSS.n7252 11.636
R11174 VSS.n7252 VSS.n7249 11.636
R11175 VSS.n7249 VSS.n7246 11.636
R11176 VSS.n7246 VSS.n7243 11.636
R11177 VSS.n7243 VSS.n7240 11.636
R11178 VSS.n7240 VSS.n7237 11.636
R11179 VSS.n7237 VSS.n7234 11.636
R11180 VSS.n7234 VSS.n7231 11.636
R11181 VSS.n7231 VSS.n7228 11.636
R11182 VSS.n7228 VSS.n7225 11.636
R11183 VSS.n9186 VSS.n9183 11.636
R11184 VSS.n9183 VSS.n9180 11.636
R11185 VSS.n9180 VSS.n9177 11.636
R11186 VSS.n9177 VSS.n9174 11.636
R11187 VSS.n9174 VSS.n9171 11.636
R11188 VSS.n9171 VSS.n9168 11.636
R11189 VSS.n9168 VSS.n9165 11.636
R11190 VSS.n9165 VSS.n9162 11.636
R11191 VSS.n9162 VSS.n9159 11.636
R11192 VSS.n9159 VSS.n9156 11.636
R11193 VSS.n9156 VSS.n9153 11.636
R11194 VSS.n8934 VSS.n8931 11.636
R11195 VSS.n8931 VSS.n8928 11.636
R11196 VSS.n8928 VSS.n8925 11.636
R11197 VSS.n8925 VSS.n8922 11.636
R11198 VSS.n8922 VSS.n8919 11.636
R11199 VSS.n8919 VSS.n8916 11.636
R11200 VSS.n8916 VSS.n8913 11.636
R11201 VSS.n8913 VSS.n8910 11.636
R11202 VSS.n8910 VSS.n8907 11.636
R11203 VSS.n9150 VSS.n9147 11.636
R11204 VSS.n8679 VSS.n8676 11.636
R11205 VSS.n8676 VSS.n8673 11.636
R11206 VSS.n8673 VSS.n8670 11.636
R11207 VSS.n8670 VSS.n8667 11.636
R11208 VSS.n8667 VSS.n8664 11.636
R11209 VSS.n8940 VSS.n8937 11.636
R11210 VSS.n8943 VSS.n8940 11.636
R11211 VSS.n8946 VSS.n8943 11.636
R11212 VSS.n8949 VSS.n8946 11.636
R11213 VSS.n8950 VSS.n8949 11.636
R11214 VSS.n8434 VSS.n8431 11.636
R11215 VSS.n8431 VSS.n8428 11.636
R11216 VSS.n8428 VSS.n8425 11.636
R11217 VSS.n8425 VSS.n8422 11.636
R11218 VSS.n8422 VSS.n8419 11.636
R11219 VSS.n8685 VSS.n8682 11.636
R11220 VSS.n8688 VSS.n8685 11.636
R11221 VSS.n8691 VSS.n8688 11.636
R11222 VSS.n8694 VSS.n8691 11.636
R11223 VSS.n8695 VSS.n8694 11.636
R11224 VSS.n8191 VSS.n8188 11.636
R11225 VSS.n8188 VSS.n8185 11.636
R11226 VSS.n8185 VSS.n8182 11.636
R11227 VSS.n8182 VSS.n8179 11.636
R11228 VSS.n8179 VSS.n8176 11.636
R11229 VSS.n8440 VSS.n8437 11.636
R11230 VSS.n8443 VSS.n8440 11.636
R11231 VSS.n8446 VSS.n8443 11.636
R11232 VSS.n8449 VSS.n8446 11.636
R11233 VSS.n8450 VSS.n8449 11.636
R11234 VSS.n7946 VSS.n7943 11.636
R11235 VSS.n7943 VSS.n7940 11.636
R11236 VSS.n7940 VSS.n7937 11.636
R11237 VSS.n7937 VSS.n7934 11.636
R11238 VSS.n7934 VSS.n7931 11.636
R11239 VSS.n8197 VSS.n8194 11.636
R11240 VSS.n8200 VSS.n8197 11.636
R11241 VSS.n8203 VSS.n8200 11.636
R11242 VSS.n8206 VSS.n8203 11.636
R11243 VSS.n8207 VSS.n8206 11.636
R11244 VSS.n7703 VSS.n7700 11.636
R11245 VSS.n7700 VSS.n7697 11.636
R11246 VSS.n7697 VSS.n7694 11.636
R11247 VSS.n7694 VSS.n7691 11.636
R11248 VSS.n7691 VSS.n7688 11.636
R11249 VSS.n7952 VSS.n7949 11.636
R11250 VSS.n7955 VSS.n7952 11.636
R11251 VSS.n7958 VSS.n7955 11.636
R11252 VSS.n7961 VSS.n7958 11.636
R11253 VSS.n7962 VSS.n7961 11.636
R11254 VSS.n7446 VSS.n7443 11.636
R11255 VSS.n7443 VSS.n7440 11.636
R11256 VSS.n7440 VSS.n7437 11.636
R11257 VSS.n7437 VSS.n7434 11.636
R11258 VSS.n7434 VSS.n7431 11.636
R11259 VSS.n7709 VSS.n7706 11.636
R11260 VSS.n7712 VSS.n7709 11.636
R11261 VSS.n7715 VSS.n7712 11.636
R11262 VSS.n7718 VSS.n7715 11.636
R11263 VSS.n7719 VSS.n7718 11.636
R11264 VSS.n7222 VSS.n7219 11.636
R11265 VSS.n7452 VSS.n7449 11.636
R11266 VSS.n7455 VSS.n7452 11.636
R11267 VSS.n7458 VSS.n7455 11.636
R11268 VSS.n7461 VSS.n7458 11.636
R11269 VSS.n7464 VSS.n7461 11.636
R11270 VSS.n7467 VSS.n7464 11.636
R11271 VSS.n7470 VSS.n7467 11.636
R11272 VSS.n7473 VSS.n7470 11.636
R11273 VSS.n7474 VSS.n7473 11.636
R11274 VSS.n1652 VSS.n1587 11.636
R11275 VSS.n1592 VSS.n1587 11.636
R11276 VSS.n1645 VSS.n1592 11.636
R11277 VSS.n1645 VSS.n1644 11.636
R11278 VSS.n1644 VSS.n1643 11.636
R11279 VSS.n1643 VSS.n1593 11.636
R11280 VSS.n1637 VSS.n1593 11.636
R11281 VSS.n1637 VSS.n1636 11.636
R11282 VSS.n1636 VSS.n1635 11.636
R11283 VSS.n1635 VSS.n1597 11.636
R11284 VSS.n1629 VSS.n1597 11.636
R11285 VSS.n1119 VSS.n637 11.636
R11286 VSS.n1119 VSS.n1115 11.636
R11287 VSS.n1125 VSS.n1115 11.636
R11288 VSS.n1126 VSS.n1125 11.636
R11289 VSS.n1127 VSS.n1126 11.636
R11290 VSS.n1127 VSS.n1111 11.636
R11291 VSS.n1133 VSS.n1111 11.636
R11292 VSS.n1134 VSS.n1133 11.636
R11293 VSS.n1135 VSS.n1134 11.636
R11294 VSS.n1135 VSS.n1107 11.636
R11295 VSS.n1141 VSS.n1107 11.636
R11296 VSS.n1165 VSS.n1095 11.636
R11297 VSS.n1159 VSS.n1095 11.636
R11298 VSS.n1159 VSS.n1158 11.636
R11299 VSS.n1158 VSS.n1157 11.636
R11300 VSS.n1157 VSS.n1099 11.636
R11301 VSS.n1151 VSS.n1099 11.636
R11302 VSS.n1151 VSS.n1150 11.636
R11303 VSS.n1150 VSS.n1149 11.636
R11304 VSS.n1149 VSS.n1103 11.636
R11305 VSS.n1143 VSS.n1103 11.636
R11306 VSS.n1143 VSS.n1142 11.636
R11307 VSS.n1321 VSS.n624 11.636
R11308 VSS.n628 VSS.n624 11.636
R11309 VSS.n1314 VSS.n628 11.636
R11310 VSS.n1314 VSS.n1313 11.636
R11311 VSS.n1313 VSS.n1312 11.636
R11312 VSS.n1312 VSS.n629 11.636
R11313 VSS.n1306 VSS.n629 11.636
R11314 VSS.n1306 VSS.n1305 11.636
R11315 VSS.n1305 VSS.n1304 11.636
R11316 VSS.n1304 VSS.n633 11.636
R11317 VSS.n1298 VSS.n633 11.636
R11318 VSS.n1348 VSS.n1347 11.636
R11319 VSS.n1347 VSS.n1346 11.636
R11320 VSS.n1346 VSS.n609 11.636
R11321 VSS.n1340 VSS.n609 11.636
R11322 VSS.n1340 VSS.n1339 11.636
R11323 VSS.n1339 VSS.n1338 11.636
R11324 VSS.n1338 VSS.n613 11.636
R11325 VSS.n1332 VSS.n613 11.636
R11326 VSS.n1332 VSS.n1331 11.636
R11327 VSS.n1331 VSS.n1330 11.636
R11328 VSS.n1330 VSS.n617 11.636
R11329 VSS.n5652 VSS.n1361 11.636
R11330 VSS.n5653 VSS.n5652 11.636
R11331 VSS.n5654 VSS.n5653 11.636
R11332 VSS.n5654 VSS.n1357 11.636
R11333 VSS.n5660 VSS.n1357 11.636
R11334 VSS.n5661 VSS.n5660 11.636
R11335 VSS.n5662 VSS.n5661 11.636
R11336 VSS.n5662 VSS.n1353 11.636
R11337 VSS.n5668 VSS.n1353 11.636
R11338 VSS.n5669 VSS.n5668 11.636
R11339 VSS.n5670 VSS.n5669 11.636
R11340 VSS.n1489 VSS.n1488 11.636
R11341 VSS.n1488 VSS.n1487 11.636
R11342 VSS.n1487 VSS.n1464 11.636
R11343 VSS.n1481 VSS.n1464 11.636
R11344 VSS.n1481 VSS.n1480 11.636
R11345 VSS.n1480 VSS.n1479 11.636
R11346 VSS.n1479 VSS.n1468 11.636
R11347 VSS.n1473 VSS.n1468 11.636
R11348 VSS.n1473 VSS.n1472 11.636
R11349 VSS.n1472 VSS.n1367 11.636
R11350 VSS.n5645 VSS.n1367 11.636
R11351 VSS.n5444 VSS.n1502 11.636
R11352 VSS.n5445 VSS.n5444 11.636
R11353 VSS.n5446 VSS.n5445 11.636
R11354 VSS.n5446 VSS.n1498 11.636
R11355 VSS.n5452 VSS.n1498 11.636
R11356 VSS.n5453 VSS.n5452 11.636
R11357 VSS.n5454 VSS.n5453 11.636
R11358 VSS.n5454 VSS.n1494 11.636
R11359 VSS.n5460 VSS.n1494 11.636
R11360 VSS.n5461 VSS.n5460 11.636
R11361 VSS.n5462 VSS.n5461 11.636
R11362 VSS.n1628 VSS.n1627 11.636
R11363 VSS.n1627 VSS.n1601 11.636
R11364 VSS.n1621 VSS.n1601 11.636
R11365 VSS.n1621 VSS.n1620 11.636
R11366 VSS.n1620 VSS.n1619 11.636
R11367 VSS.n1619 VSS.n1605 11.636
R11368 VSS.n1613 VSS.n1605 11.636
R11369 VSS.n1613 VSS.n1612 11.636
R11370 VSS.n1612 VSS.n1611 11.636
R11371 VSS.n1611 VSS.n1508 11.636
R11372 VSS.n5437 VSS.n1508 11.636
R11373 VSS.n3815 VSS.n3814 11.636
R11374 VSS.n3816 VSS.n3815 11.636
R11375 VSS.n3816 VSS.n3442 11.636
R11376 VSS.n3822 VSS.n3442 11.636
R11377 VSS.n3823 VSS.n3822 11.636
R11378 VSS.n3824 VSS.n3823 11.636
R11379 VSS.n3824 VSS.n3438 11.636
R11380 VSS.n3830 VSS.n3438 11.636
R11381 VSS.n3831 VSS.n3830 11.636
R11382 VSS.n3832 VSS.n3831 11.636
R11383 VSS.n3832 VSS.n3434 11.636
R11384 VSS.n5128 VSS.n3097 11.636
R11385 VSS.n5122 VSS.n3097 11.636
R11386 VSS.n5122 VSS.n5121 11.636
R11387 VSS.n5121 VSS.n5120 11.636
R11388 VSS.n5120 VSS.n3103 11.636
R11389 VSS.n5114 VSS.n3103 11.636
R11390 VSS.n5114 VSS.n5113 11.636
R11391 VSS.n5113 VSS.n5112 11.636
R11392 VSS.n5112 VSS.n3107 11.636
R11393 VSS.n5106 VSS.n3107 11.636
R11394 VSS.n5106 VSS.n5105 11.636
R11395 VSS.n5082 VSS.n5081 11.636
R11396 VSS.n5082 VSS.n3119 11.636
R11397 VSS.n5088 VSS.n3119 11.636
R11398 VSS.n5089 VSS.n5088 11.636
R11399 VSS.n5090 VSS.n5089 11.636
R11400 VSS.n5090 VSS.n3115 11.636
R11401 VSS.n5096 VSS.n3115 11.636
R11402 VSS.n5097 VSS.n5096 11.636
R11403 VSS.n5098 VSS.n5097 11.636
R11404 VSS.n5098 VSS.n3111 11.636
R11405 VSS.n5104 VSS.n3111 11.636
R11406 VSS.n5054 VSS.n5053 11.636
R11407 VSS.n5055 VSS.n5054 11.636
R11408 VSS.n5055 VSS.n3134 11.636
R11409 VSS.n5061 VSS.n3134 11.636
R11410 VSS.n5062 VSS.n5061 11.636
R11411 VSS.n5063 VSS.n5062 11.636
R11412 VSS.n5063 VSS.n3130 11.636
R11413 VSS.n5070 VSS.n3130 11.636
R11414 VSS.n5071 VSS.n5070 11.636
R11415 VSS.n5072 VSS.n5071 11.636
R11416 VSS.n5072 VSS.n3123 11.636
R11417 VSS.n3275 VSS.n3274 11.636
R11418 VSS.n3274 VSS.n3273 11.636
R11419 VSS.n3273 VSS.n3245 11.636
R11420 VSS.n3267 VSS.n3245 11.636
R11421 VSS.n3267 VSS.n3266 11.636
R11422 VSS.n3266 VSS.n3265 11.636
R11423 VSS.n3265 VSS.n3249 11.636
R11424 VSS.n3259 VSS.n3249 11.636
R11425 VSS.n3259 VSS.n3258 11.636
R11426 VSS.n3258 VSS.n3257 11.636
R11427 VSS.n3257 VSS.n3253 11.636
R11428 VSS.n4482 VSS.n3288 11.636
R11429 VSS.n4483 VSS.n4482 11.636
R11430 VSS.n4484 VSS.n4483 11.636
R11431 VSS.n4484 VSS.n3284 11.636
R11432 VSS.n4490 VSS.n3284 11.636
R11433 VSS.n4491 VSS.n4490 11.636
R11434 VSS.n4492 VSS.n4491 11.636
R11435 VSS.n4492 VSS.n3280 11.636
R11436 VSS.n4498 VSS.n3280 11.636
R11437 VSS.n4499 VSS.n4498 11.636
R11438 VSS.n4500 VSS.n4499 11.636
R11439 VSS.n4449 VSS.n3303 11.636
R11440 VSS.n4455 VSS.n3303 11.636
R11441 VSS.n4456 VSS.n4455 11.636
R11442 VSS.n4457 VSS.n4456 11.636
R11443 VSS.n4457 VSS.n3299 11.636
R11444 VSS.n4463 VSS.n3299 11.636
R11445 VSS.n4464 VSS.n4463 11.636
R11446 VSS.n4466 VSS.n4464 11.636
R11447 VSS.n4466 VSS.n4465 11.636
R11448 VSS.n4465 VSS.n3295 11.636
R11449 VSS.n4473 VSS.n3295 11.636
R11450 VSS.n3917 VSS.n3405 11.636
R11451 VSS.n3917 VSS.n3916 11.636
R11452 VSS.n3916 VSS.n3915 11.636
R11453 VSS.n3915 VSS.n3889 11.636
R11454 VSS.n3909 VSS.n3889 11.636
R11455 VSS.n3909 VSS.n3908 11.636
R11456 VSS.n3908 VSS.n3907 11.636
R11457 VSS.n3907 VSS.n3894 11.636
R11458 VSS.n3901 VSS.n3894 11.636
R11459 VSS.n3901 VSS.n3900 11.636
R11460 VSS.n3900 VSS.n3307 11.636
R11461 VSS.n3867 VSS.n3866 11.636
R11462 VSS.n3867 VSS.n3415 11.636
R11463 VSS.n3873 VSS.n3415 11.636
R11464 VSS.n3874 VSS.n3873 11.636
R11465 VSS.n3875 VSS.n3874 11.636
R11466 VSS.n3875 VSS.n3411 11.636
R11467 VSS.n3881 VSS.n3411 11.636
R11468 VSS.n3882 VSS.n3881 11.636
R11469 VSS.n3883 VSS.n3882 11.636
R11470 VSS.n3883 VSS.n3406 11.636
R11471 VSS.n3924 VSS.n3406 11.636
R11472 VSS.n3839 VSS.n3838 11.636
R11473 VSS.n3840 VSS.n3839 11.636
R11474 VSS.n3840 VSS.n3430 11.636
R11475 VSS.n3846 VSS.n3430 11.636
R11476 VSS.n3847 VSS.n3846 11.636
R11477 VSS.n3848 VSS.n3847 11.636
R11478 VSS.n3848 VSS.n3426 11.636
R11479 VSS.n3855 VSS.n3426 11.636
R11480 VSS.n3856 VSS.n3855 11.636
R11481 VSS.n3857 VSS.n3856 11.636
R11482 VSS.n3857 VSS.n3419 11.636
R11483 VSS.n17849 VSS.n17809 11.636
R11484 VSS.n17849 VSS.n17848 11.636
R11485 VSS.n17848 VSS.n17847 11.636
R11486 VSS.n17847 VSS.n17811 11.636
R11487 VSS.n17841 VSS.n17811 11.636
R11488 VSS.n17841 VSS.n17840 11.636
R11489 VSS.n17840 VSS.n17839 11.636
R11490 VSS.n17839 VSS.n17816 11.636
R11491 VSS.n17833 VSS.n17816 11.636
R11492 VSS.n17833 VSS.n17832 11.636
R11493 VSS.n17832 VSS.n17831 11.636
R11494 VSS.n17857 VSS.n17856 11.636
R11495 VSS.n17858 VSS.n17857 11.636
R11496 VSS.n17858 VSS.n17801 11.636
R11497 VSS.n17864 VSS.n17801 11.636
R11498 VSS.n17865 VSS.n17864 11.636
R11499 VSS.n17866 VSS.n17865 11.636
R11500 VSS.n17872 VSS.n17797 11.636
R11501 VSS.n17873 VSS.n17872 11.636
R11502 VSS.n17874 VSS.n17873 11.636
R11503 VSS.n17874 VSS.n17793 11.636
R11504 VSS.n17882 VSS.n17881 11.636
R11505 VSS.n17882 VSS.n17789 11.636
R11506 VSS.n17888 VSS.n17789 11.636
R11507 VSS.n17889 VSS.n17888 11.636
R11508 VSS.n17890 VSS.n17889 11.636
R11509 VSS.n17890 VSS.n17785 11.636
R11510 VSS.n17896 VSS.n17785 11.636
R11511 VSS.n17897 VSS.n17896 11.636
R11512 VSS.n17898 VSS.n17897 11.636
R11513 VSS.n17898 VSS.n17781 11.636
R11514 VSS.n17904 VSS.n17781 11.636
R11515 VSS.n17825 VSS.n17820 11.636
R11516 VSS.n17825 VSS.n17824 11.636
R11517 VSS.n17824 VSS.n17770 11.636
R11518 VSS.n17920 VSS.n17771 11.636
R11519 VSS.n17914 VSS.n17771 11.636
R11520 VSS.n17914 VSS.n17913 11.636
R11521 VSS.n17913 VSS.n17912 11.636
R11522 VSS.n17912 VSS.n17777 11.636
R11523 VSS.n17906 VSS.n17777 11.636
R11524 VSS.n17906 VSS.n17905 11.636
R11525 VSS VSS.n10578 10.944
R11526 VSS VSS.n18230 10.83
R11527 VSS.n17610 VSS.n17598 10.438
R11528 VSS VSS.n17797 10.343
R11529 VSS.n2455 VSS.n2324 9.955
R11530 VSS.n2448 VSS.n2447 9.955
R11531 VSS.n2387 VSS.n2384 9.955
R11532 VSS.n2435 VSS.n2390 9.955
R11533 VSS.n2429 VSS.n2394 9.955
R11534 VSS.n2423 VSS.n2397 9.955
R11535 VSS.n2418 VSS.n2400 9.955
R11536 VSS.n2412 VSS.n2403 9.955
R11537 VSS.n2545 VSS.n2234 9.955
R11538 VSS.n2538 VSS.n2537 9.955
R11539 VSS.n2477 VSS.n2474 9.955
R11540 VSS.n2525 VSS.n2480 9.955
R11541 VSS.n2519 VSS.n2484 9.955
R11542 VSS.n2513 VSS.n2487 9.955
R11543 VSS.n2508 VSS.n2490 9.955
R11544 VSS.n2502 VSS.n2493 9.955
R11545 VSS.n2635 VSS.n2144 9.955
R11546 VSS.n2628 VSS.n2627 9.955
R11547 VSS.n2567 VSS.n2564 9.955
R11548 VSS.n2615 VSS.n2570 9.955
R11549 VSS.n2609 VSS.n2574 9.955
R11550 VSS.n2603 VSS.n2577 9.955
R11551 VSS.n2598 VSS.n2580 9.955
R11552 VSS.n2592 VSS.n2583 9.955
R11553 VSS.n2725 VSS.n2054 9.955
R11554 VSS.n2718 VSS.n2717 9.955
R11555 VSS.n2657 VSS.n2654 9.955
R11556 VSS.n2705 VSS.n2660 9.955
R11557 VSS.n2699 VSS.n2664 9.955
R11558 VSS.n2693 VSS.n2667 9.955
R11559 VSS.n2688 VSS.n2670 9.955
R11560 VSS.n2682 VSS.n2673 9.955
R11561 VSS.n2815 VSS.n1964 9.955
R11562 VSS.n2808 VSS.n2807 9.955
R11563 VSS.n2747 VSS.n2744 9.955
R11564 VSS.n2795 VSS.n2750 9.955
R11565 VSS.n2789 VSS.n2754 9.955
R11566 VSS.n2783 VSS.n2757 9.955
R11567 VSS.n2778 VSS.n2760 9.955
R11568 VSS.n2772 VSS.n2763 9.955
R11569 VSS.n2905 VSS.n1874 9.955
R11570 VSS.n2898 VSS.n2897 9.955
R11571 VSS.n2837 VSS.n2834 9.955
R11572 VSS.n2885 VSS.n2840 9.955
R11573 VSS.n2879 VSS.n2844 9.955
R11574 VSS.n2873 VSS.n2847 9.955
R11575 VSS.n2868 VSS.n2850 9.955
R11576 VSS.n2862 VSS.n2853 9.955
R11577 VSS.n2995 VSS.n1784 9.955
R11578 VSS.n2988 VSS.n2987 9.955
R11579 VSS.n2927 VSS.n2924 9.955
R11580 VSS.n2975 VSS.n2930 9.955
R11581 VSS.n2969 VSS.n2934 9.955
R11582 VSS.n2963 VSS.n2937 9.955
R11583 VSS.n2958 VSS.n2940 9.955
R11584 VSS.n2952 VSS.n2943 9.955
R11585 VSS.n3085 VSS.n1694 9.955
R11586 VSS.n3078 VSS.n3077 9.955
R11587 VSS.n3017 VSS.n3014 9.955
R11588 VSS.n3065 VSS.n3020 9.955
R11589 VSS.n3059 VSS.n3024 9.955
R11590 VSS.n3053 VSS.n3027 9.955
R11591 VSS.n3048 VSS.n3030 9.955
R11592 VSS.n3042 VSS.n3033 9.955
R11593 VSS.n6131 VSS.n6130 9.955
R11594 VSS.n6139 VSS.n6138 9.955
R11595 VSS.n6147 VSS.n6146 9.955
R11596 VSS.n6155 VSS.n6154 9.955
R11597 VSS.n6163 VSS.n6162 9.955
R11598 VSS.n6171 VSS.n6170 9.955
R11599 VSS.n6179 VSS.n6178 9.955
R11600 VSS.n6187 VSS.n6186 9.955
R11601 VSS.n6015 VSS.n6014 9.955
R11602 VSS.n6023 VSS.n6022 9.955
R11603 VSS.n6031 VSS.n6030 9.955
R11604 VSS.n6039 VSS.n6038 9.955
R11605 VSS.n6047 VSS.n6046 9.955
R11606 VSS.n6055 VSS.n6054 9.955
R11607 VSS.n6063 VSS.n6062 9.955
R11608 VSS.n6071 VSS.n6070 9.955
R11609 VSS.n5899 VSS.n5898 9.955
R11610 VSS.n5907 VSS.n5906 9.955
R11611 VSS.n5915 VSS.n5914 9.955
R11612 VSS.n5923 VSS.n5922 9.955
R11613 VSS.n5931 VSS.n5930 9.955
R11614 VSS.n5939 VSS.n5938 9.955
R11615 VSS.n5947 VSS.n5946 9.955
R11616 VSS.n5955 VSS.n5954 9.955
R11617 VSS.n7039 VSS.n5791 9.955
R11618 VSS.n7033 VSS.n5796 9.955
R11619 VSS.n7027 VSS.n5802 9.955
R11620 VSS.n7021 VSS.n5808 9.955
R11621 VSS.n7015 VSS.n5814 9.955
R11622 VSS.n7009 VSS.n5819 9.955
R11623 VSS.n7003 VSS.n5826 9.955
R11624 VSS.n6997 VSS.n5832 9.955
R11625 VSS.n6928 VSS.n6438 9.955
R11626 VSS.n6921 VSS.n6920 9.955
R11627 VSS.n6861 VSS.n6858 9.955
R11628 VSS.n6908 VSS.n6864 9.955
R11629 VSS.n6902 VSS.n6868 9.955
R11630 VSS.n6896 VSS.n6872 9.955
R11631 VSS.n6890 VSS.n6875 9.955
R11632 VSS.n6885 VSS.n6878 9.955
R11633 VSS.n6838 VSS.n6528 9.955
R11634 VSS.n6831 VSS.n6830 9.955
R11635 VSS.n6771 VSS.n6768 9.955
R11636 VSS.n6818 VSS.n6774 9.955
R11637 VSS.n6812 VSS.n6778 9.955
R11638 VSS.n6806 VSS.n6782 9.955
R11639 VSS.n6800 VSS.n6785 9.955
R11640 VSS.n6795 VSS.n6788 9.955
R11641 VSS.n6748 VSS.n6618 9.955
R11642 VSS.n6741 VSS.n6740 9.955
R11643 VSS.n6681 VSS.n6678 9.955
R11644 VSS.n6728 VSS.n6684 9.955
R11645 VSS.n6722 VSS.n6688 9.955
R11646 VSS.n6716 VSS.n6692 9.955
R11647 VSS.n6710 VSS.n6695 9.955
R11648 VSS.n6705 VSS.n6698 9.955
R11649 VSS.n16522 VSS.n16521 9.3
R11650 VSS.n16521 VSS.n16520 9.3
R11651 VSS.n16508 VSS.n16507 9.3
R11652 VSS.n16507 VSS.n16506 9.3
R11653 VSS.n16494 VSS.n16493 9.3
R11654 VSS.n16493 VSS.n16492 9.3
R11655 VSS.n16480 VSS.n16479 9.3
R11656 VSS.n16479 VSS.n16478 9.3
R11657 VSS.n16471 VSS.n16470 9.3
R11658 VSS.n16473 VSS.n16471 9.3
R11659 VSS.n16473 VSS.n16472 9.3
R11660 VSS.n16462 VSS.n16461 9.3
R11661 VSS.n16461 VSS.n16460 9.3
R11662 VSS.n16444 VSS.n16443 9.3
R11663 VSS.n16443 VSS.n16442 9.3
R11664 VSS.n16430 VSS.n16429 9.3
R11665 VSS.n16429 VSS.n16428 9.3
R11666 VSS.n16416 VSS.n16415 9.3
R11667 VSS.n16415 VSS.n16414 9.3
R11668 VSS.n16402 VSS.n16401 9.3
R11669 VSS.n16401 VSS.n16400 9.3
R11670 VSS.n16388 VSS.n16387 9.3
R11671 VSS.n16387 VSS.n16386 9.3
R11672 VSS.n16284 VSS.n16283 9.3
R11673 VSS.n16283 VSS.n16282 9.3
R11674 VSS.n16266 VSS.n16265 9.3
R11675 VSS.n16265 VSS.n16264 9.3
R11676 VSS.n16252 VSS.n16251 9.3
R11677 VSS.n16251 VSS.n16250 9.3
R11678 VSS.n16238 VSS.n16237 9.3
R11679 VSS.n16237 VSS.n16236 9.3
R11680 VSS.n16224 VSS.n16223 9.3
R11681 VSS.n16223 VSS.n16222 9.3
R11682 VSS.n16215 VSS.n16214 9.3
R11683 VSS.n16217 VSS.n16215 9.3
R11684 VSS.n16217 VSS.n16216 9.3
R11685 VSS.n16206 VSS.n16205 9.3
R11686 VSS.n16205 VSS.n16204 9.3
R11687 VSS.n16188 VSS.n16187 9.3
R11688 VSS.n16187 VSS.n16186 9.3
R11689 VSS.n16174 VSS.n16173 9.3
R11690 VSS.n16173 VSS.n16172 9.3
R11691 VSS.n16160 VSS.n16159 9.3
R11692 VSS.n16159 VSS.n16158 9.3
R11693 VSS.n16146 VSS.n16145 9.3
R11694 VSS.n16145 VSS.n16144 9.3
R11695 VSS.n16132 VSS.n16131 9.3
R11696 VSS.n16131 VSS.n16130 9.3
R11697 VSS.n16040 VSS.n16039 9.3
R11698 VSS.n16039 VSS.n16038 9.3
R11699 VSS.n16022 VSS.n16021 9.3
R11700 VSS.n16021 VSS.n16020 9.3
R11701 VSS.n16008 VSS.n16007 9.3
R11702 VSS.n16007 VSS.n16006 9.3
R11703 VSS.n15994 VSS.n15993 9.3
R11704 VSS.n15993 VSS.n15992 9.3
R11705 VSS.n15980 VSS.n15979 9.3
R11706 VSS.n15979 VSS.n15978 9.3
R11707 VSS.n15971 VSS.n15970 9.3
R11708 VSS.n15973 VSS.n15971 9.3
R11709 VSS.n15973 VSS.n15972 9.3
R11710 VSS.n15962 VSS.n15961 9.3
R11711 VSS.n15961 VSS.n15960 9.3
R11712 VSS.n15944 VSS.n15943 9.3
R11713 VSS.n15943 VSS.n15942 9.3
R11714 VSS.n15930 VSS.n15929 9.3
R11715 VSS.n15929 VSS.n15928 9.3
R11716 VSS.n15916 VSS.n15915 9.3
R11717 VSS.n15915 VSS.n15914 9.3
R11718 VSS.n15902 VSS.n15901 9.3
R11719 VSS.n15901 VSS.n15900 9.3
R11720 VSS.n15888 VSS.n15887 9.3
R11721 VSS.n15887 VSS.n15886 9.3
R11722 VSS.n15796 VSS.n15795 9.3
R11723 VSS.n15795 VSS.n15794 9.3
R11724 VSS.n15778 VSS.n15777 9.3
R11725 VSS.n15777 VSS.n15776 9.3
R11726 VSS.n15764 VSS.n15763 9.3
R11727 VSS.n15763 VSS.n15762 9.3
R11728 VSS.n15750 VSS.n15749 9.3
R11729 VSS.n15749 VSS.n15748 9.3
R11730 VSS.n15736 VSS.n15735 9.3
R11731 VSS.n15735 VSS.n15734 9.3
R11732 VSS.n15727 VSS.n15726 9.3
R11733 VSS.n15729 VSS.n15727 9.3
R11734 VSS.n15729 VSS.n15728 9.3
R11735 VSS.n15718 VSS.n15717 9.3
R11736 VSS.n15717 VSS.n15716 9.3
R11737 VSS.n15700 VSS.n15699 9.3
R11738 VSS.n15699 VSS.n15698 9.3
R11739 VSS.n15686 VSS.n15685 9.3
R11740 VSS.n15685 VSS.n15684 9.3
R11741 VSS.n15672 VSS.n15671 9.3
R11742 VSS.n15671 VSS.n15670 9.3
R11743 VSS.n15658 VSS.n15657 9.3
R11744 VSS.n15657 VSS.n15656 9.3
R11745 VSS.n15644 VSS.n15643 9.3
R11746 VSS.n15643 VSS.n15642 9.3
R11747 VSS.n15552 VSS.n15551 9.3
R11748 VSS.n15551 VSS.n15550 9.3
R11749 VSS.n15534 VSS.n15533 9.3
R11750 VSS.n15533 VSS.n15532 9.3
R11751 VSS.n15520 VSS.n15519 9.3
R11752 VSS.n15519 VSS.n15518 9.3
R11753 VSS.n15506 VSS.n15505 9.3
R11754 VSS.n15505 VSS.n15504 9.3
R11755 VSS.n15492 VSS.n15491 9.3
R11756 VSS.n15491 VSS.n15490 9.3
R11757 VSS.n15483 VSS.n15482 9.3
R11758 VSS.n15485 VSS.n15483 9.3
R11759 VSS.n15485 VSS.n15484 9.3
R11760 VSS.n15474 VSS.n15473 9.3
R11761 VSS.n15473 VSS.n15472 9.3
R11762 VSS.n15456 VSS.n15455 9.3
R11763 VSS.n15455 VSS.n15454 9.3
R11764 VSS.n15442 VSS.n15441 9.3
R11765 VSS.n15441 VSS.n15440 9.3
R11766 VSS.n15428 VSS.n15427 9.3
R11767 VSS.n15427 VSS.n15426 9.3
R11768 VSS.n15414 VSS.n15413 9.3
R11769 VSS.n15413 VSS.n15412 9.3
R11770 VSS.n15400 VSS.n15399 9.3
R11771 VSS.n15399 VSS.n15398 9.3
R11772 VSS.n15308 VSS.n15307 9.3
R11773 VSS.n15307 VSS.n15306 9.3
R11774 VSS.n15290 VSS.n15289 9.3
R11775 VSS.n15289 VSS.n15288 9.3
R11776 VSS.n15276 VSS.n15275 9.3
R11777 VSS.n15275 VSS.n15274 9.3
R11778 VSS.n15262 VSS.n15261 9.3
R11779 VSS.n15261 VSS.n15260 9.3
R11780 VSS.n15248 VSS.n15247 9.3
R11781 VSS.n15247 VSS.n15246 9.3
R11782 VSS.n15239 VSS.n15238 9.3
R11783 VSS.n15241 VSS.n15239 9.3
R11784 VSS.n15241 VSS.n15240 9.3
R11785 VSS.n15230 VSS.n15229 9.3
R11786 VSS.n15229 VSS.n15228 9.3
R11787 VSS.n15212 VSS.n15211 9.3
R11788 VSS.n15211 VSS.n15210 9.3
R11789 VSS.n15198 VSS.n15197 9.3
R11790 VSS.n15197 VSS.n15196 9.3
R11791 VSS.n15184 VSS.n15183 9.3
R11792 VSS.n15183 VSS.n15182 9.3
R11793 VSS.n15170 VSS.n15169 9.3
R11794 VSS.n15169 VSS.n15168 9.3
R11795 VSS.n15156 VSS.n15155 9.3
R11796 VSS.n15155 VSS.n15154 9.3
R11797 VSS.n15064 VSS.n15063 9.3
R11798 VSS.n15063 VSS.n15062 9.3
R11799 VSS.n15046 VSS.n15045 9.3
R11800 VSS.n15045 VSS.n15044 9.3
R11801 VSS.n15032 VSS.n15031 9.3
R11802 VSS.n15031 VSS.n15030 9.3
R11803 VSS.n15018 VSS.n15017 9.3
R11804 VSS.n15017 VSS.n15016 9.3
R11805 VSS.n15004 VSS.n15003 9.3
R11806 VSS.n15003 VSS.n15002 9.3
R11807 VSS.n14995 VSS.n14994 9.3
R11808 VSS.n14997 VSS.n14995 9.3
R11809 VSS.n14997 VSS.n14996 9.3
R11810 VSS.n14986 VSS.n14985 9.3
R11811 VSS.n14985 VSS.n14984 9.3
R11812 VSS.n14968 VSS.n14967 9.3
R11813 VSS.n14967 VSS.n14966 9.3
R11814 VSS.n14954 VSS.n14953 9.3
R11815 VSS.n14953 VSS.n14952 9.3
R11816 VSS.n14940 VSS.n14939 9.3
R11817 VSS.n14939 VSS.n14938 9.3
R11818 VSS.n14926 VSS.n14925 9.3
R11819 VSS.n14925 VSS.n14924 9.3
R11820 VSS.n14912 VSS.n14911 9.3
R11821 VSS.n14911 VSS.n14910 9.3
R11822 VSS.n14808 VSS.n14807 9.3
R11823 VSS.n14807 VSS.n14806 9.3
R11824 VSS.n14790 VSS.n14789 9.3
R11825 VSS.n14789 VSS.n14788 9.3
R11826 VSS.n14776 VSS.n14775 9.3
R11827 VSS.n14775 VSS.n14774 9.3
R11828 VSS.n14762 VSS.n14761 9.3
R11829 VSS.n14761 VSS.n14760 9.3
R11830 VSS.n14748 VSS.n14747 9.3
R11831 VSS.n14747 VSS.n14746 9.3
R11832 VSS.n14739 VSS.n14738 9.3
R11833 VSS.n14741 VSS.n14739 9.3
R11834 VSS.n14741 VSS.n14740 9.3
R11835 VSS.n14730 VSS.n14729 9.3
R11836 VSS.n14729 VSS.n14728 9.3
R11837 VSS.n14712 VSS.n14711 9.3
R11838 VSS.n14711 VSS.n14710 9.3
R11839 VSS.n14698 VSS.n14697 9.3
R11840 VSS.n14697 VSS.n14696 9.3
R11841 VSS.n14684 VSS.n14683 9.3
R11842 VSS.n14683 VSS.n14682 9.3
R11843 VSS.n14670 VSS.n14669 9.3
R11844 VSS.n14669 VSS.n14668 9.3
R11845 VSS.n14656 VSS.n14655 9.3
R11846 VSS.n14655 VSS.n14654 9.3
R11847 VSS.n16583 VSS.n16582 9.3
R11848 VSS.n16582 VSS.n16581 9.3
R11849 VSS.n16598 VSS.n16597 9.3
R11850 VSS.n16610 VSS.n16609 9.3
R11851 VSS.n16622 VSS.n16621 9.3
R11852 VSS.n16638 VSS.n16637 9.3
R11853 VSS.n16637 VSS.n16636 9.3
R11854 VSS.n16646 VSS.n16645 9.3
R11855 VSS.n16658 VSS.n16657 9.3
R11856 VSS.n16670 VSS.n16669 9.3
R11857 VSS.n16682 VSS.n16681 9.3
R11858 VSS.n16741 VSS.n16740 9.3
R11859 VSS.n16766 VSS.n16765 9.3
R11860 VSS.n16778 VSS.n16777 9.3
R11861 VSS.n16790 VSS.n16789 9.3
R11862 VSS.n16806 VSS.n16805 9.3
R11863 VSS.n16805 VSS.n16804 9.3
R11864 VSS.n16814 VSS.n16813 9.3
R11865 VSS.n16826 VSS.n16825 9.3
R11866 VSS.n16838 VSS.n16837 9.3
R11867 VSS.n16850 VSS.n16849 9.3
R11868 VSS.n16909 VSS.n16908 9.3
R11869 VSS.n16934 VSS.n16933 9.3
R11870 VSS.n16946 VSS.n16945 9.3
R11871 VSS.n16958 VSS.n16957 9.3
R11872 VSS.n16974 VSS.n16973 9.3
R11873 VSS.n16973 VSS.n16972 9.3
R11874 VSS.n16982 VSS.n16981 9.3
R11875 VSS.n16994 VSS.n16993 9.3
R11876 VSS.n17006 VSS.n17005 9.3
R11877 VSS.n17018 VSS.n17017 9.3
R11878 VSS.n17077 VSS.n17076 9.3
R11879 VSS.n17102 VSS.n17101 9.3
R11880 VSS.n17114 VSS.n17113 9.3
R11881 VSS.n17126 VSS.n17125 9.3
R11882 VSS.n17142 VSS.n17141 9.3
R11883 VSS.n17141 VSS.n17140 9.3
R11884 VSS.n17150 VSS.n17149 9.3
R11885 VSS.n17162 VSS.n17161 9.3
R11886 VSS.n17174 VSS.n17173 9.3
R11887 VSS.n17186 VSS.n17185 9.3
R11888 VSS.n17245 VSS.n17244 9.3
R11889 VSS.n17270 VSS.n17269 9.3
R11890 VSS.n17282 VSS.n17281 9.3
R11891 VSS.n17294 VSS.n17293 9.3
R11892 VSS.n17310 VSS.n17309 9.3
R11893 VSS.n17309 VSS.n17308 9.3
R11894 VSS.n17318 VSS.n17317 9.3
R11895 VSS.n17330 VSS.n17329 9.3
R11896 VSS.n17342 VSS.n17341 9.3
R11897 VSS.n17354 VSS.n17353 9.3
R11898 VSS.n17413 VSS.n17412 9.3
R11899 VSS.n17438 VSS.n17437 9.3
R11900 VSS.n17450 VSS.n17449 9.3
R11901 VSS.n17462 VSS.n17461 9.3
R11902 VSS.n17478 VSS.n17477 9.3
R11903 VSS.n17477 VSS.n17476 9.3
R11904 VSS.n17486 VSS.n17485 9.3
R11905 VSS.n17498 VSS.n17497 9.3
R11906 VSS.n17510 VSS.n17509 9.3
R11907 VSS.n17522 VSS.n17521 9.3
R11908 VSS.n17581 VSS.n17580 9.3
R11909 VSS.n14224 VSS.n14223 9.3
R11910 VSS.n14212 VSS.n14211 9.3
R11911 VSS.n14200 VSS.n14193 9.3
R11912 VSS.n14200 VSS.n14199 9.3
R11913 VSS.n14188 VSS.n14187 9.3
R11914 VSS.n14176 VSS.n14175 9.3
R11915 VSS.n14164 VSS.n14163 9.3
R11916 VSS.n14152 VSS.n14151 9.3
R11917 VSS.n14140 VSS.n14139 9.3
R11918 VSS.n14281 VSS.n14280 9.3
R11919 VSS.n14404 VSS.n14403 9.3
R11920 VSS.n14392 VSS.n14391 9.3
R11921 VSS.n14380 VSS.n14373 9.3
R11922 VSS.n14380 VSS.n14379 9.3
R11923 VSS.n14368 VSS.n14367 9.3
R11924 VSS.n14356 VSS.n14355 9.3
R11925 VSS.n14344 VSS.n14343 9.3
R11926 VSS.n14332 VSS.n14331 9.3
R11927 VSS.n14320 VSS.n14319 9.3
R11928 VSS.n14461 VSS.n14460 9.3
R11929 VSS.n12571 VSS.n12570 9.3
R11930 VSS.n12570 VSS.n12569 9.3
R11931 VSS.n12557 VSS.n12556 9.3
R11932 VSS.n12556 VSS.n12555 9.3
R11933 VSS.n12543 VSS.n12542 9.3
R11934 VSS.n12542 VSS.n12541 9.3
R11935 VSS.n12529 VSS.n12528 9.3
R11936 VSS.n12528 VSS.n12527 9.3
R11937 VSS.n12520 VSS.n12519 9.3
R11938 VSS.n12522 VSS.n12520 9.3
R11939 VSS.n12522 VSS.n12521 9.3
R11940 VSS.n12511 VSS.n12510 9.3
R11941 VSS.n12510 VSS.n12509 9.3
R11942 VSS.n12493 VSS.n12492 9.3
R11943 VSS.n12492 VSS.n12491 9.3
R11944 VSS.n12479 VSS.n12478 9.3
R11945 VSS.n12478 VSS.n12477 9.3
R11946 VSS.n12465 VSS.n12464 9.3
R11947 VSS.n12464 VSS.n12463 9.3
R11948 VSS.n12451 VSS.n12450 9.3
R11949 VSS.n12450 VSS.n12449 9.3
R11950 VSS.n12437 VSS.n12436 9.3
R11951 VSS.n12436 VSS.n12435 9.3
R11952 VSS.n12333 VSS.n12332 9.3
R11953 VSS.n12332 VSS.n12331 9.3
R11954 VSS.n12315 VSS.n12314 9.3
R11955 VSS.n12314 VSS.n12313 9.3
R11956 VSS.n12301 VSS.n12300 9.3
R11957 VSS.n12300 VSS.n12299 9.3
R11958 VSS.n12287 VSS.n12286 9.3
R11959 VSS.n12286 VSS.n12285 9.3
R11960 VSS.n12273 VSS.n12272 9.3
R11961 VSS.n12272 VSS.n12271 9.3
R11962 VSS.n12264 VSS.n12263 9.3
R11963 VSS.n12266 VSS.n12264 9.3
R11964 VSS.n12266 VSS.n12265 9.3
R11965 VSS.n12255 VSS.n12254 9.3
R11966 VSS.n12254 VSS.n12253 9.3
R11967 VSS.n12237 VSS.n12236 9.3
R11968 VSS.n12236 VSS.n12235 9.3
R11969 VSS.n12223 VSS.n12222 9.3
R11970 VSS.n12222 VSS.n12221 9.3
R11971 VSS.n12209 VSS.n12208 9.3
R11972 VSS.n12208 VSS.n12207 9.3
R11973 VSS.n12195 VSS.n12194 9.3
R11974 VSS.n12194 VSS.n12193 9.3
R11975 VSS.n12181 VSS.n12180 9.3
R11976 VSS.n12180 VSS.n12179 9.3
R11977 VSS.n12089 VSS.n12088 9.3
R11978 VSS.n12088 VSS.n12087 9.3
R11979 VSS.n12071 VSS.n12070 9.3
R11980 VSS.n12070 VSS.n12069 9.3
R11981 VSS.n12057 VSS.n12056 9.3
R11982 VSS.n12056 VSS.n12055 9.3
R11983 VSS.n12043 VSS.n12042 9.3
R11984 VSS.n12042 VSS.n12041 9.3
R11985 VSS.n12029 VSS.n12028 9.3
R11986 VSS.n12028 VSS.n12027 9.3
R11987 VSS.n12020 VSS.n12019 9.3
R11988 VSS.n12022 VSS.n12020 9.3
R11989 VSS.n12022 VSS.n12021 9.3
R11990 VSS.n12011 VSS.n12010 9.3
R11991 VSS.n12010 VSS.n12009 9.3
R11992 VSS.n11993 VSS.n11992 9.3
R11993 VSS.n11992 VSS.n11991 9.3
R11994 VSS.n11979 VSS.n11978 9.3
R11995 VSS.n11978 VSS.n11977 9.3
R11996 VSS.n11965 VSS.n11964 9.3
R11997 VSS.n11964 VSS.n11963 9.3
R11998 VSS.n11951 VSS.n11950 9.3
R11999 VSS.n11950 VSS.n11949 9.3
R12000 VSS.n11937 VSS.n11936 9.3
R12001 VSS.n11936 VSS.n11935 9.3
R12002 VSS.n11845 VSS.n11844 9.3
R12003 VSS.n11844 VSS.n11843 9.3
R12004 VSS.n11827 VSS.n11826 9.3
R12005 VSS.n11826 VSS.n11825 9.3
R12006 VSS.n11813 VSS.n11812 9.3
R12007 VSS.n11812 VSS.n11811 9.3
R12008 VSS.n11799 VSS.n11798 9.3
R12009 VSS.n11798 VSS.n11797 9.3
R12010 VSS.n11785 VSS.n11784 9.3
R12011 VSS.n11784 VSS.n11783 9.3
R12012 VSS.n11776 VSS.n11775 9.3
R12013 VSS.n11778 VSS.n11776 9.3
R12014 VSS.n11778 VSS.n11777 9.3
R12015 VSS.n11767 VSS.n11766 9.3
R12016 VSS.n11766 VSS.n11765 9.3
R12017 VSS.n11749 VSS.n11748 9.3
R12018 VSS.n11748 VSS.n11747 9.3
R12019 VSS.n11735 VSS.n11734 9.3
R12020 VSS.n11734 VSS.n11733 9.3
R12021 VSS.n11721 VSS.n11720 9.3
R12022 VSS.n11720 VSS.n11719 9.3
R12023 VSS.n11707 VSS.n11706 9.3
R12024 VSS.n11706 VSS.n11705 9.3
R12025 VSS.n11693 VSS.n11692 9.3
R12026 VSS.n11692 VSS.n11691 9.3
R12027 VSS.n11601 VSS.n11600 9.3
R12028 VSS.n11600 VSS.n11599 9.3
R12029 VSS.n11583 VSS.n11582 9.3
R12030 VSS.n11582 VSS.n11581 9.3
R12031 VSS.n11569 VSS.n11568 9.3
R12032 VSS.n11568 VSS.n11567 9.3
R12033 VSS.n11555 VSS.n11554 9.3
R12034 VSS.n11554 VSS.n11553 9.3
R12035 VSS.n11541 VSS.n11540 9.3
R12036 VSS.n11540 VSS.n11539 9.3
R12037 VSS.n11532 VSS.n11531 9.3
R12038 VSS.n11534 VSS.n11532 9.3
R12039 VSS.n11534 VSS.n11533 9.3
R12040 VSS.n11523 VSS.n11522 9.3
R12041 VSS.n11522 VSS.n11521 9.3
R12042 VSS.n11505 VSS.n11504 9.3
R12043 VSS.n11504 VSS.n11503 9.3
R12044 VSS.n11491 VSS.n11490 9.3
R12045 VSS.n11490 VSS.n11489 9.3
R12046 VSS.n11477 VSS.n11476 9.3
R12047 VSS.n11476 VSS.n11475 9.3
R12048 VSS.n11463 VSS.n11462 9.3
R12049 VSS.n11462 VSS.n11461 9.3
R12050 VSS.n11449 VSS.n11448 9.3
R12051 VSS.n11448 VSS.n11447 9.3
R12052 VSS.n11357 VSS.n11356 9.3
R12053 VSS.n11356 VSS.n11355 9.3
R12054 VSS.n11339 VSS.n11338 9.3
R12055 VSS.n11338 VSS.n11337 9.3
R12056 VSS.n11325 VSS.n11324 9.3
R12057 VSS.n11324 VSS.n11323 9.3
R12058 VSS.n11311 VSS.n11310 9.3
R12059 VSS.n11310 VSS.n11309 9.3
R12060 VSS.n11297 VSS.n11296 9.3
R12061 VSS.n11296 VSS.n11295 9.3
R12062 VSS.n11288 VSS.n11287 9.3
R12063 VSS.n11290 VSS.n11288 9.3
R12064 VSS.n11290 VSS.n11289 9.3
R12065 VSS.n11279 VSS.n11278 9.3
R12066 VSS.n11278 VSS.n11277 9.3
R12067 VSS.n11261 VSS.n11260 9.3
R12068 VSS.n11260 VSS.n11259 9.3
R12069 VSS.n11247 VSS.n11246 9.3
R12070 VSS.n11246 VSS.n11245 9.3
R12071 VSS.n11233 VSS.n11232 9.3
R12072 VSS.n11232 VSS.n11231 9.3
R12073 VSS.n11219 VSS.n11218 9.3
R12074 VSS.n11218 VSS.n11217 9.3
R12075 VSS.n11205 VSS.n11204 9.3
R12076 VSS.n11204 VSS.n11203 9.3
R12077 VSS.n11113 VSS.n11112 9.3
R12078 VSS.n11112 VSS.n11111 9.3
R12079 VSS.n11095 VSS.n11094 9.3
R12080 VSS.n11094 VSS.n11093 9.3
R12081 VSS.n11081 VSS.n11080 9.3
R12082 VSS.n11080 VSS.n11079 9.3
R12083 VSS.n11067 VSS.n11066 9.3
R12084 VSS.n11066 VSS.n11065 9.3
R12085 VSS.n11053 VSS.n11052 9.3
R12086 VSS.n11052 VSS.n11051 9.3
R12087 VSS.n11044 VSS.n11043 9.3
R12088 VSS.n11046 VSS.n11044 9.3
R12089 VSS.n11046 VSS.n11045 9.3
R12090 VSS.n11035 VSS.n11034 9.3
R12091 VSS.n11034 VSS.n11033 9.3
R12092 VSS.n11017 VSS.n11016 9.3
R12093 VSS.n11016 VSS.n11015 9.3
R12094 VSS.n11003 VSS.n11002 9.3
R12095 VSS.n11002 VSS.n11001 9.3
R12096 VSS.n10989 VSS.n10988 9.3
R12097 VSS.n10988 VSS.n10987 9.3
R12098 VSS.n10975 VSS.n10974 9.3
R12099 VSS.n10974 VSS.n10973 9.3
R12100 VSS.n10961 VSS.n10960 9.3
R12101 VSS.n10960 VSS.n10959 9.3
R12102 VSS.n10857 VSS.n10856 9.3
R12103 VSS.n10856 VSS.n10855 9.3
R12104 VSS.n10839 VSS.n10838 9.3
R12105 VSS.n10838 VSS.n10837 9.3
R12106 VSS.n10825 VSS.n10824 9.3
R12107 VSS.n10824 VSS.n10823 9.3
R12108 VSS.n10811 VSS.n10810 9.3
R12109 VSS.n10810 VSS.n10809 9.3
R12110 VSS.n10797 VSS.n10796 9.3
R12111 VSS.n10796 VSS.n10795 9.3
R12112 VSS.n10788 VSS.n10787 9.3
R12113 VSS.n10790 VSS.n10788 9.3
R12114 VSS.n10790 VSS.n10789 9.3
R12115 VSS.n10779 VSS.n10778 9.3
R12116 VSS.n10778 VSS.n10777 9.3
R12117 VSS.n10761 VSS.n10760 9.3
R12118 VSS.n10760 VSS.n10759 9.3
R12119 VSS.n10747 VSS.n10746 9.3
R12120 VSS.n10746 VSS.n10745 9.3
R12121 VSS.n10733 VSS.n10732 9.3
R12122 VSS.n10732 VSS.n10731 9.3
R12123 VSS.n10719 VSS.n10718 9.3
R12124 VSS.n10718 VSS.n10717 9.3
R12125 VSS.n10705 VSS.n10704 9.3
R12126 VSS.n10704 VSS.n10703 9.3
R12127 VSS.n12632 VSS.n12631 9.3
R12128 VSS.n12631 VSS.n12630 9.3
R12129 VSS.n12741 VSS.n12740 9.3
R12130 VSS.n12729 VSS.n12728 9.3
R12131 VSS.n12717 VSS.n12710 9.3
R12132 VSS.n12717 VSS.n12716 9.3
R12133 VSS.n12705 VSS.n12704 9.3
R12134 VSS.n12693 VSS.n12692 9.3
R12135 VSS.n12681 VSS.n12680 9.3
R12136 VSS.n12669 VSS.n12668 9.3
R12137 VSS.n12657 VSS.n12656 9.3
R12138 VSS.n12798 VSS.n12797 9.3
R12139 VSS.n12921 VSS.n12920 9.3
R12140 VSS.n12909 VSS.n12908 9.3
R12141 VSS.n12897 VSS.n12890 9.3
R12142 VSS.n12897 VSS.n12896 9.3
R12143 VSS.n12885 VSS.n12884 9.3
R12144 VSS.n12873 VSS.n12872 9.3
R12145 VSS.n12861 VSS.n12860 9.3
R12146 VSS.n12849 VSS.n12848 9.3
R12147 VSS.n12837 VSS.n12836 9.3
R12148 VSS.n12978 VSS.n12977 9.3
R12149 VSS.n13101 VSS.n13100 9.3
R12150 VSS.n13089 VSS.n13088 9.3
R12151 VSS.n13077 VSS.n13070 9.3
R12152 VSS.n13077 VSS.n13076 9.3
R12153 VSS.n13065 VSS.n13064 9.3
R12154 VSS.n13053 VSS.n13052 9.3
R12155 VSS.n13041 VSS.n13040 9.3
R12156 VSS.n13029 VSS.n13028 9.3
R12157 VSS.n13017 VSS.n13016 9.3
R12158 VSS.n13158 VSS.n13157 9.3
R12159 VSS.n13281 VSS.n13280 9.3
R12160 VSS.n13269 VSS.n13268 9.3
R12161 VSS.n13257 VSS.n13250 9.3
R12162 VSS.n13257 VSS.n13256 9.3
R12163 VSS.n13245 VSS.n13244 9.3
R12164 VSS.n13233 VSS.n13232 9.3
R12165 VSS.n13221 VSS.n13220 9.3
R12166 VSS.n13209 VSS.n13208 9.3
R12167 VSS.n13197 VSS.n13196 9.3
R12168 VSS.n13338 VSS.n13337 9.3
R12169 VSS.n13461 VSS.n13460 9.3
R12170 VSS.n13449 VSS.n13448 9.3
R12171 VSS.n13437 VSS.n13430 9.3
R12172 VSS.n13437 VSS.n13436 9.3
R12173 VSS.n13425 VSS.n13424 9.3
R12174 VSS.n13413 VSS.n13412 9.3
R12175 VSS.n13401 VSS.n13400 9.3
R12176 VSS.n13389 VSS.n13388 9.3
R12177 VSS.n13377 VSS.n13376 9.3
R12178 VSS.n13518 VSS.n13517 9.3
R12179 VSS.n13641 VSS.n13640 9.3
R12180 VSS.n13629 VSS.n13628 9.3
R12181 VSS.n13617 VSS.n13610 9.3
R12182 VSS.n13617 VSS.n13616 9.3
R12183 VSS.n13605 VSS.n13604 9.3
R12184 VSS.n13593 VSS.n13592 9.3
R12185 VSS.n13581 VSS.n13580 9.3
R12186 VSS.n13569 VSS.n13568 9.3
R12187 VSS.n13557 VSS.n13556 9.3
R12188 VSS.n13698 VSS.n13697 9.3
R12189 VSS.n13821 VSS.n13820 9.3
R12190 VSS.n13809 VSS.n13808 9.3
R12191 VSS.n13797 VSS.n13790 9.3
R12192 VSS.n13797 VSS.n13796 9.3
R12193 VSS.n13785 VSS.n13784 9.3
R12194 VSS.n13773 VSS.n13772 9.3
R12195 VSS.n13761 VSS.n13760 9.3
R12196 VSS.n13749 VSS.n13748 9.3
R12197 VSS.n13737 VSS.n13736 9.3
R12198 VSS.n13878 VSS.n13877 9.3
R12199 VSS.n14001 VSS.n14000 9.3
R12200 VSS.n13989 VSS.n13988 9.3
R12201 VSS.n13977 VSS.n13970 9.3
R12202 VSS.n13977 VSS.n13976 9.3
R12203 VSS.n13965 VSS.n13964 9.3
R12204 VSS.n13953 VSS.n13952 9.3
R12205 VSS.n13941 VSS.n13940 9.3
R12206 VSS.n13929 VSS.n13928 9.3
R12207 VSS.n13917 VSS.n13916 9.3
R12208 VSS.n14058 VSS.n14057 9.3
R12209 VSS.n9139 VSS.n9138 9.3
R12210 VSS.n9138 VSS.n9137 9.3
R12211 VSS.n9125 VSS.n9124 9.3
R12212 VSS.n9124 VSS.n9123 9.3
R12213 VSS.n9111 VSS.n9110 9.3
R12214 VSS.n9110 VSS.n9109 9.3
R12215 VSS.n9097 VSS.n9096 9.3
R12216 VSS.n9096 VSS.n9095 9.3
R12217 VSS.n9088 VSS.n9087 9.3
R12218 VSS.n9090 VSS.n9088 9.3
R12219 VSS.n9090 VSS.n9089 9.3
R12220 VSS.n9079 VSS.n9078 9.3
R12221 VSS.n9078 VSS.n9077 9.3
R12222 VSS.n9061 VSS.n9060 9.3
R12223 VSS.n9060 VSS.n9059 9.3
R12224 VSS.n9047 VSS.n9046 9.3
R12225 VSS.n9046 VSS.n9045 9.3
R12226 VSS.n9033 VSS.n9032 9.3
R12227 VSS.n9032 VSS.n9031 9.3
R12228 VSS.n9019 VSS.n9018 9.3
R12229 VSS.n9018 VSS.n9017 9.3
R12230 VSS.n9005 VSS.n9004 9.3
R12231 VSS.n9004 VSS.n9003 9.3
R12232 VSS.n8901 VSS.n8900 9.3
R12233 VSS.n8900 VSS.n8899 9.3
R12234 VSS.n8883 VSS.n8882 9.3
R12235 VSS.n8882 VSS.n8881 9.3
R12236 VSS.n8869 VSS.n8868 9.3
R12237 VSS.n8868 VSS.n8867 9.3
R12238 VSS.n8855 VSS.n8854 9.3
R12239 VSS.n8854 VSS.n8853 9.3
R12240 VSS.n8841 VSS.n8840 9.3
R12241 VSS.n8840 VSS.n8839 9.3
R12242 VSS.n8832 VSS.n8831 9.3
R12243 VSS.n8834 VSS.n8832 9.3
R12244 VSS.n8834 VSS.n8833 9.3
R12245 VSS.n8823 VSS.n8822 9.3
R12246 VSS.n8822 VSS.n8821 9.3
R12247 VSS.n8805 VSS.n8804 9.3
R12248 VSS.n8804 VSS.n8803 9.3
R12249 VSS.n8791 VSS.n8790 9.3
R12250 VSS.n8790 VSS.n8789 9.3
R12251 VSS.n8777 VSS.n8776 9.3
R12252 VSS.n8776 VSS.n8775 9.3
R12253 VSS.n8763 VSS.n8762 9.3
R12254 VSS.n8762 VSS.n8761 9.3
R12255 VSS.n8749 VSS.n8748 9.3
R12256 VSS.n8748 VSS.n8747 9.3
R12257 VSS.n8657 VSS.n8656 9.3
R12258 VSS.n8656 VSS.n8655 9.3
R12259 VSS.n8639 VSS.n8638 9.3
R12260 VSS.n8638 VSS.n8637 9.3
R12261 VSS.n8625 VSS.n8624 9.3
R12262 VSS.n8624 VSS.n8623 9.3
R12263 VSS.n8611 VSS.n8610 9.3
R12264 VSS.n8610 VSS.n8609 9.3
R12265 VSS.n8597 VSS.n8596 9.3
R12266 VSS.n8596 VSS.n8595 9.3
R12267 VSS.n8588 VSS.n8587 9.3
R12268 VSS.n8590 VSS.n8588 9.3
R12269 VSS.n8590 VSS.n8589 9.3
R12270 VSS.n8579 VSS.n8578 9.3
R12271 VSS.n8578 VSS.n8577 9.3
R12272 VSS.n8561 VSS.n8560 9.3
R12273 VSS.n8560 VSS.n8559 9.3
R12274 VSS.n8547 VSS.n8546 9.3
R12275 VSS.n8546 VSS.n8545 9.3
R12276 VSS.n8533 VSS.n8532 9.3
R12277 VSS.n8532 VSS.n8531 9.3
R12278 VSS.n8519 VSS.n8518 9.3
R12279 VSS.n8518 VSS.n8517 9.3
R12280 VSS.n8505 VSS.n8504 9.3
R12281 VSS.n8504 VSS.n8503 9.3
R12282 VSS.n8413 VSS.n8412 9.3
R12283 VSS.n8412 VSS.n8411 9.3
R12284 VSS.n8395 VSS.n8394 9.3
R12285 VSS.n8394 VSS.n8393 9.3
R12286 VSS.n8381 VSS.n8380 9.3
R12287 VSS.n8380 VSS.n8379 9.3
R12288 VSS.n8367 VSS.n8366 9.3
R12289 VSS.n8366 VSS.n8365 9.3
R12290 VSS.n8353 VSS.n8352 9.3
R12291 VSS.n8352 VSS.n8351 9.3
R12292 VSS.n8344 VSS.n8343 9.3
R12293 VSS.n8346 VSS.n8344 9.3
R12294 VSS.n8346 VSS.n8345 9.3
R12295 VSS.n8335 VSS.n8334 9.3
R12296 VSS.n8334 VSS.n8333 9.3
R12297 VSS.n8317 VSS.n8316 9.3
R12298 VSS.n8316 VSS.n8315 9.3
R12299 VSS.n8303 VSS.n8302 9.3
R12300 VSS.n8302 VSS.n8301 9.3
R12301 VSS.n8289 VSS.n8288 9.3
R12302 VSS.n8288 VSS.n8287 9.3
R12303 VSS.n8275 VSS.n8274 9.3
R12304 VSS.n8274 VSS.n8273 9.3
R12305 VSS.n8261 VSS.n8260 9.3
R12306 VSS.n8260 VSS.n8259 9.3
R12307 VSS.n8169 VSS.n8168 9.3
R12308 VSS.n8168 VSS.n8167 9.3
R12309 VSS.n8151 VSS.n8150 9.3
R12310 VSS.n8150 VSS.n8149 9.3
R12311 VSS.n8137 VSS.n8136 9.3
R12312 VSS.n8136 VSS.n8135 9.3
R12313 VSS.n8123 VSS.n8122 9.3
R12314 VSS.n8122 VSS.n8121 9.3
R12315 VSS.n8109 VSS.n8108 9.3
R12316 VSS.n8108 VSS.n8107 9.3
R12317 VSS.n8100 VSS.n8099 9.3
R12318 VSS.n8102 VSS.n8100 9.3
R12319 VSS.n8102 VSS.n8101 9.3
R12320 VSS.n8091 VSS.n8090 9.3
R12321 VSS.n8090 VSS.n8089 9.3
R12322 VSS.n8073 VSS.n8072 9.3
R12323 VSS.n8072 VSS.n8071 9.3
R12324 VSS.n8059 VSS.n8058 9.3
R12325 VSS.n8058 VSS.n8057 9.3
R12326 VSS.n8045 VSS.n8044 9.3
R12327 VSS.n8044 VSS.n8043 9.3
R12328 VSS.n8031 VSS.n8030 9.3
R12329 VSS.n8030 VSS.n8029 9.3
R12330 VSS.n8017 VSS.n8016 9.3
R12331 VSS.n8016 VSS.n8015 9.3
R12332 VSS.n7925 VSS.n7924 9.3
R12333 VSS.n7924 VSS.n7923 9.3
R12334 VSS.n7907 VSS.n7906 9.3
R12335 VSS.n7906 VSS.n7905 9.3
R12336 VSS.n7893 VSS.n7892 9.3
R12337 VSS.n7892 VSS.n7891 9.3
R12338 VSS.n7879 VSS.n7878 9.3
R12339 VSS.n7878 VSS.n7877 9.3
R12340 VSS.n7865 VSS.n7864 9.3
R12341 VSS.n7864 VSS.n7863 9.3
R12342 VSS.n7856 VSS.n7855 9.3
R12343 VSS.n7858 VSS.n7856 9.3
R12344 VSS.n7858 VSS.n7857 9.3
R12345 VSS.n7847 VSS.n7846 9.3
R12346 VSS.n7846 VSS.n7845 9.3
R12347 VSS.n7829 VSS.n7828 9.3
R12348 VSS.n7828 VSS.n7827 9.3
R12349 VSS.n7815 VSS.n7814 9.3
R12350 VSS.n7814 VSS.n7813 9.3
R12351 VSS.n7801 VSS.n7800 9.3
R12352 VSS.n7800 VSS.n7799 9.3
R12353 VSS.n7787 VSS.n7786 9.3
R12354 VSS.n7786 VSS.n7785 9.3
R12355 VSS.n7773 VSS.n7772 9.3
R12356 VSS.n7772 VSS.n7771 9.3
R12357 VSS.n7681 VSS.n7680 9.3
R12358 VSS.n7680 VSS.n7679 9.3
R12359 VSS.n7663 VSS.n7662 9.3
R12360 VSS.n7662 VSS.n7661 9.3
R12361 VSS.n7649 VSS.n7648 9.3
R12362 VSS.n7648 VSS.n7647 9.3
R12363 VSS.n7635 VSS.n7634 9.3
R12364 VSS.n7634 VSS.n7633 9.3
R12365 VSS.n7621 VSS.n7620 9.3
R12366 VSS.n7620 VSS.n7619 9.3
R12367 VSS.n7612 VSS.n7611 9.3
R12368 VSS.n7614 VSS.n7612 9.3
R12369 VSS.n7614 VSS.n7613 9.3
R12370 VSS.n7603 VSS.n7602 9.3
R12371 VSS.n7602 VSS.n7601 9.3
R12372 VSS.n7585 VSS.n7584 9.3
R12373 VSS.n7584 VSS.n7583 9.3
R12374 VSS.n7571 VSS.n7570 9.3
R12375 VSS.n7570 VSS.n7569 9.3
R12376 VSS.n7557 VSS.n7556 9.3
R12377 VSS.n7556 VSS.n7555 9.3
R12378 VSS.n7543 VSS.n7542 9.3
R12379 VSS.n7542 VSS.n7541 9.3
R12380 VSS.n7529 VSS.n7528 9.3
R12381 VSS.n7528 VSS.n7527 9.3
R12382 VSS.n7425 VSS.n7424 9.3
R12383 VSS.n7424 VSS.n7423 9.3
R12384 VSS.n7407 VSS.n7406 9.3
R12385 VSS.n7406 VSS.n7405 9.3
R12386 VSS.n7393 VSS.n7392 9.3
R12387 VSS.n7392 VSS.n7391 9.3
R12388 VSS.n7379 VSS.n7378 9.3
R12389 VSS.n7378 VSS.n7377 9.3
R12390 VSS.n7365 VSS.n7364 9.3
R12391 VSS.n7364 VSS.n7363 9.3
R12392 VSS.n7356 VSS.n7355 9.3
R12393 VSS.n7358 VSS.n7356 9.3
R12394 VSS.n7358 VSS.n7357 9.3
R12395 VSS.n7347 VSS.n7346 9.3
R12396 VSS.n7346 VSS.n7345 9.3
R12397 VSS.n7329 VSS.n7328 9.3
R12398 VSS.n7328 VSS.n7327 9.3
R12399 VSS.n7315 VSS.n7314 9.3
R12400 VSS.n7314 VSS.n7313 9.3
R12401 VSS.n7301 VSS.n7300 9.3
R12402 VSS.n7300 VSS.n7299 9.3
R12403 VSS.n7287 VSS.n7286 9.3
R12404 VSS.n7286 VSS.n7285 9.3
R12405 VSS.n7273 VSS.n7272 9.3
R12406 VSS.n7272 VSS.n7271 9.3
R12407 VSS.n9200 VSS.n9199 9.3
R12408 VSS.n9199 VSS.n9198 9.3
R12409 VSS.n10248 VSS.n10247 9.3
R12410 VSS.n10260 VSS.n10259 9.3
R12411 VSS.n10276 VSS.n10275 9.3
R12412 VSS.n10275 VSS.n10274 9.3
R12413 VSS.n10284 VSS.n10283 9.3
R12414 VSS.n10296 VSS.n10295 9.3
R12415 VSS.n10308 VSS.n10307 9.3
R12416 VSS.n10320 VSS.n10319 9.3
R12417 VSS.n10377 VSS.n10376 9.3
R12418 VSS.n10236 VSS.n10235 9.3
R12419 VSS.n10080 VSS.n10079 9.3
R12420 VSS.n10092 VSS.n10091 9.3
R12421 VSS.n10108 VSS.n10107 9.3
R12422 VSS.n10107 VSS.n10106 9.3
R12423 VSS.n10116 VSS.n10115 9.3
R12424 VSS.n10128 VSS.n10127 9.3
R12425 VSS.n10140 VSS.n10139 9.3
R12426 VSS.n10152 VSS.n10151 9.3
R12427 VSS.n10209 VSS.n10208 9.3
R12428 VSS.n10068 VSS.n10067 9.3
R12429 VSS.n9912 VSS.n9911 9.3
R12430 VSS.n9924 VSS.n9923 9.3
R12431 VSS.n9940 VSS.n9939 9.3
R12432 VSS.n9939 VSS.n9938 9.3
R12433 VSS.n9948 VSS.n9947 9.3
R12434 VSS.n9960 VSS.n9959 9.3
R12435 VSS.n9972 VSS.n9971 9.3
R12436 VSS.n9984 VSS.n9983 9.3
R12437 VSS.n10041 VSS.n10040 9.3
R12438 VSS.n9900 VSS.n9899 9.3
R12439 VSS.n9744 VSS.n9743 9.3
R12440 VSS.n9756 VSS.n9755 9.3
R12441 VSS.n9772 VSS.n9771 9.3
R12442 VSS.n9771 VSS.n9770 9.3
R12443 VSS.n9780 VSS.n9779 9.3
R12444 VSS.n9792 VSS.n9791 9.3
R12445 VSS.n9804 VSS.n9803 9.3
R12446 VSS.n9816 VSS.n9815 9.3
R12447 VSS.n9873 VSS.n9872 9.3
R12448 VSS.n9732 VSS.n9731 9.3
R12449 VSS.n9576 VSS.n9575 9.3
R12450 VSS.n9588 VSS.n9587 9.3
R12451 VSS.n9604 VSS.n9603 9.3
R12452 VSS.n9603 VSS.n9602 9.3
R12453 VSS.n9612 VSS.n9611 9.3
R12454 VSS.n9624 VSS.n9623 9.3
R12455 VSS.n9636 VSS.n9635 9.3
R12456 VSS.n9648 VSS.n9647 9.3
R12457 VSS.n9705 VSS.n9704 9.3
R12458 VSS.n9564 VSS.n9563 9.3
R12459 VSS.n9408 VSS.n9407 9.3
R12460 VSS.n9420 VSS.n9419 9.3
R12461 VSS.n9436 VSS.n9435 9.3
R12462 VSS.n9435 VSS.n9434 9.3
R12463 VSS.n9444 VSS.n9443 9.3
R12464 VSS.n9456 VSS.n9455 9.3
R12465 VSS.n9468 VSS.n9467 9.3
R12466 VSS.n9480 VSS.n9479 9.3
R12467 VSS.n9537 VSS.n9536 9.3
R12468 VSS.n9396 VSS.n9395 9.3
R12469 VSS.n9240 VSS.n9239 9.3
R12470 VSS.n9252 VSS.n9251 9.3
R12471 VSS.n9268 VSS.n9267 9.3
R12472 VSS.n9267 VSS.n9266 9.3
R12473 VSS.n9276 VSS.n9275 9.3
R12474 VSS.n9288 VSS.n9287 9.3
R12475 VSS.n9300 VSS.n9299 9.3
R12476 VSS.n9312 VSS.n9311 9.3
R12477 VSS.n9369 VSS.n9368 9.3
R12478 VSS.n9228 VSS.n9227 9.3
R12479 VSS.n10403 VSS.n10402 9.3
R12480 VSS.n10427 VSS.n10426 9.3
R12481 VSS.n10451 VSS.n10450 9.3
R12482 VSS.n10475 VSS.n10474 9.3
R12483 VSS.n10545 VSS.n10544 9.3
R12484 VSS.n10487 VSS.n10486 9.3
R12485 VSS.n10463 VSS.n10462 9.3
R12486 VSS.n10443 VSS.n10442 9.3
R12487 VSS.n10442 VSS.n10441 9.3
R12488 VSS.n10415 VSS.n10414 9.3
R12489 VSS.n4850 VSS.n4849 9.3
R12490 VSS.n4850 VSS.n4828 9.3
R12491 VSS.n4828 VSS.n4827 9.3
R12492 VSS.n4832 VSS.n4831 9.3
R12493 VSS.n4858 VSS.n4857 9.3
R12494 VSS.n4857 VSS.n4856 9.3
R12495 VSS.n4856 VSS.n4855 9.3
R12496 VSS.n4862 VSS.n4814 9.3
R12497 VSS.n4863 VSS.n4862 9.3
R12498 VSS.n4864 VSS.n4863 9.3
R12499 VSS.n4870 VSS.n4869 9.3
R12500 VSS.n4873 VSS.n4872 9.3
R12501 VSS.n4873 VSS.n4809 9.3
R12502 VSS.n4809 VSS.n4808 9.3
R12503 VSS.n4881 VSS.n4880 9.3
R12504 VSS.n4880 VSS.n4879 9.3
R12505 VSS.n4879 VSS.n4878 9.3
R12506 VSS.n4882 VSS.n4800 9.3
R12507 VSS.n4885 VSS.n4795 9.3
R12508 VSS.n4886 VSS.n4885 9.3
R12509 VSS.n4887 VSS.n4886 9.3
R12510 VSS.n4896 VSS.n4895 9.3
R12511 VSS.n4896 VSS.n4790 9.3
R12512 VSS.n4790 VSS.n4789 9.3
R12513 VSS.n4794 VSS.n4793 9.3
R12514 VSS.n4904 VSS.n4903 9.3
R12515 VSS.n4903 VSS.n4902 9.3
R12516 VSS.n4902 VSS.n4901 9.3
R12517 VSS.n4908 VSS.n4776 9.3
R12518 VSS.n4909 VSS.n4908 9.3
R12519 VSS.n4910 VSS.n4909 9.3
R12520 VSS.n4916 VSS.n4915 9.3
R12521 VSS.n4919 VSS.n4918 9.3
R12522 VSS.n4919 VSS.n4771 9.3
R12523 VSS.n4771 VSS.n4770 9.3
R12524 VSS.n4927 VSS.n4926 9.3
R12525 VSS.n4926 VSS.n4925 9.3
R12526 VSS.n4925 VSS.n4924 9.3
R12527 VSS.n4847 VSS.n4846 9.3
R12528 VSS.n4859 VSS.n4819 9.3
R12529 VSS.n4813 VSS.n4812 9.3
R12530 VSS.n4893 VSS.n4892 9.3
R12531 VSS.n4905 VSS.n4781 9.3
R12532 VSS.n4775 VSS.n4774 9.3
R12533 VSS.n4929 VSS.n4726 9.3
R12534 VSS.n4932 VSS.n4721 9.3
R12535 VSS.n4933 VSS.n4932 9.3
R12536 VSS.n4934 VSS.n4933 9.3
R12537 VSS.n4940 VSS.n4939 9.3
R12538 VSS.n4943 VSS.n4942 9.3
R12539 VSS.n4943 VSS.n4716 9.3
R12540 VSS.n4716 VSS.n4715 9.3
R12541 VSS.n4720 VSS.n4719 9.3
R12542 VSS.n4951 VSS.n4950 9.3
R12543 VSS.n4950 VSS.n4949 9.3
R12544 VSS.n4949 VSS.n4948 9.3
R12545 VSS.n4952 VSS.n4707 9.3
R12546 VSS.n4955 VSS.n4702 9.3
R12547 VSS.n4956 VSS.n4955 9.3
R12548 VSS.n4957 VSS.n4956 9.3
R12549 VSS.n4963 VSS.n4962 9.3
R12550 VSS.n4966 VSS.n4965 9.3
R12551 VSS.n4966 VSS.n4697 9.3
R12552 VSS.n4697 VSS.n4696 9.3
R12553 VSS.n4701 VSS.n4700 9.3
R12554 VSS.n4974 VSS.n4973 9.3
R12555 VSS.n4973 VSS.n4972 9.3
R12556 VSS.n4972 VSS.n4971 9.3
R12557 VSS.n4975 VSS.n4688 9.3
R12558 VSS.n4978 VSS.n4683 9.3
R12559 VSS.n4979 VSS.n4978 9.3
R12560 VSS.n4980 VSS.n4979 9.3
R12561 VSS.n4986 VSS.n4985 9.3
R12562 VSS.n4989 VSS.n4988 9.3
R12563 VSS.n4989 VSS.n4678 9.3
R12564 VSS.n4678 VSS.n4677 9.3
R12565 VSS.n4682 VSS.n4681 9.3
R12566 VSS.n4997 VSS.n4996 9.3
R12567 VSS.n4996 VSS.n4995 9.3
R12568 VSS.n4995 VSS.n4994 9.3
R12569 VSS.n4998 VSS.n4669 9.3
R12570 VSS.n5001 VSS.n4664 9.3
R12571 VSS.n5002 VSS.n5001 9.3
R12572 VSS.n5003 VSS.n5002 9.3
R12573 VSS.n5009 VSS.n5008 9.3
R12574 VSS.n5012 VSS.n5011 9.3
R12575 VSS.n5012 VSS.n4659 9.3
R12576 VSS.n4659 VSS.n4658 9.3
R12577 VSS.n4663 VSS.n4662 9.3
R12578 VSS.n5020 VSS.n5019 9.3
R12579 VSS.n5019 VSS.n5018 9.3
R12580 VSS.n5018 VSS.n5017 9.3
R12581 VSS.n4649 VSS.n3156 9.3
R12582 VSS.n4646 VSS.n3157 9.3
R12583 VSS.n4646 VSS.n4645 9.3
R12584 VSS.n4645 VSS.n4644 9.3
R12585 VSS.n4639 VSS.n4638 9.3
R12586 VSS.n4636 VSS.n4635 9.3
R12587 VSS.n4635 VSS.n3161 9.3
R12588 VSS.n3161 VSS.n3160 9.3
R12589 VSS.n3169 VSS.n3163 9.3
R12590 VSS.n4628 VSS.n4627 9.3
R12591 VSS.n4629 VSS.n4628 9.3
R12592 VSS.n4630 VSS.n4629 9.3
R12593 VSS.n4625 VSS.n4624 9.3
R12594 VSS.n4616 VSS.n4615 9.3
R12595 VSS.n4616 VSS.n3173 9.3
R12596 VSS.n4620 VSS.n3173 9.3
R12597 VSS.n4614 VSS.n4613 9.3
R12598 VSS.n4611 VSS.n3179 9.3
R12599 VSS.n4611 VSS.n4610 9.3
R12600 VSS.n4610 VSS.n4609 9.3
R12601 VSS.n4604 VSS.n4603 9.3
R12602 VSS.n4601 VSS.n4600 9.3
R12603 VSS.n4600 VSS.n3182 9.3
R12604 VSS.n3182 VSS.n3181 9.3
R12605 VSS.n3190 VSS.n3184 9.3
R12606 VSS.n4593 VSS.n4592 9.3
R12607 VSS.n4594 VSS.n4593 9.3
R12608 VSS.n4595 VSS.n4594 9.3
R12609 VSS.n4590 VSS.n4589 9.3
R12610 VSS.n4581 VSS.n4580 9.3
R12611 VSS.n4581 VSS.n3194 9.3
R12612 VSS.n4585 VSS.n3194 9.3
R12613 VSS.n4579 VSS.n4578 9.3
R12614 VSS.n4576 VSS.n3200 9.3
R12615 VSS.n4576 VSS.n4575 9.3
R12616 VSS.n4575 VSS.n4574 9.3
R12617 VSS.n4569 VSS.n4568 9.3
R12618 VSS.n4566 VSS.n4565 9.3
R12619 VSS.n4565 VSS.n3203 9.3
R12620 VSS.n3203 VSS.n3202 9.3
R12621 VSS.n3211 VSS.n3205 9.3
R12622 VSS.n4558 VSS.n4557 9.3
R12623 VSS.n4559 VSS.n4558 9.3
R12624 VSS.n4560 VSS.n4559 9.3
R12625 VSS.n4555 VSS.n4554 9.3
R12626 VSS.n4546 VSS.n4545 9.3
R12627 VSS.n4546 VSS.n3215 9.3
R12628 VSS.n4550 VSS.n3215 9.3
R12629 VSS.n4542 VSS.n3219 9.3
R12630 VSS.n4539 VSS.n3221 9.3
R12631 VSS.n4531 VSS.n3221 9.3
R12632 VSS.n4532 VSS.n4531 9.3
R12633 VSS.n4538 VSS.n4537 9.3
R12634 VSS.n4241 VSS.n4240 9.3
R12635 VSS.n4241 VSS.n3225 9.3
R12636 VSS.n3227 VSS.n3225 9.3
R12637 VSS.n4239 VSS.n4238 9.3
R12638 VSS.n4249 VSS.n4248 9.3
R12639 VSS.n4248 VSS.n4247 9.3
R12640 VSS.n4247 VSS.n4246 9.3
R12641 VSS.n4250 VSS.n4229 9.3
R12642 VSS.n4253 VSS.n4224 9.3
R12643 VSS.n4254 VSS.n4253 9.3
R12644 VSS.n4255 VSS.n4254 9.3
R12645 VSS.n4261 VSS.n4260 9.3
R12646 VSS.n4264 VSS.n4263 9.3
R12647 VSS.n4264 VSS.n4219 9.3
R12648 VSS.n4219 VSS.n4218 9.3
R12649 VSS.n4223 VSS.n4222 9.3
R12650 VSS.n4272 VSS.n4271 9.3
R12651 VSS.n4271 VSS.n4270 9.3
R12652 VSS.n4270 VSS.n4269 9.3
R12653 VSS.n4273 VSS.n4210 9.3
R12654 VSS.n4276 VSS.n4205 9.3
R12655 VSS.n4277 VSS.n4276 9.3
R12656 VSS.n4278 VSS.n4277 9.3
R12657 VSS.n4284 VSS.n4283 9.3
R12658 VSS.n4287 VSS.n4286 9.3
R12659 VSS.n4287 VSS.n4200 9.3
R12660 VSS.n4200 VSS.n4199 9.3
R12661 VSS.n4204 VSS.n4203 9.3
R12662 VSS.n4295 VSS.n4294 9.3
R12663 VSS.n4294 VSS.n4293 9.3
R12664 VSS.n4293 VSS.n4292 9.3
R12665 VSS.n4296 VSS.n4191 9.3
R12666 VSS.n4299 VSS.n4186 9.3
R12667 VSS.n4300 VSS.n4299 9.3
R12668 VSS.n4301 VSS.n4300 9.3
R12669 VSS.n4307 VSS.n4306 9.3
R12670 VSS.n4310 VSS.n4309 9.3
R12671 VSS.n4310 VSS.n4181 9.3
R12672 VSS.n4181 VSS.n4180 9.3
R12673 VSS.n4185 VSS.n4184 9.3
R12674 VSS.n4318 VSS.n4317 9.3
R12675 VSS.n4317 VSS.n4316 9.3
R12676 VSS.n4316 VSS.n4315 9.3
R12677 VSS.n4320 VSS.n4136 9.3
R12678 VSS.n4323 VSS.n4131 9.3
R12679 VSS.n4324 VSS.n4323 9.3
R12680 VSS.n4325 VSS.n4324 9.3
R12681 VSS.n4331 VSS.n4330 9.3
R12682 VSS.n4334 VSS.n4333 9.3
R12683 VSS.n4334 VSS.n4126 9.3
R12684 VSS.n4126 VSS.n4125 9.3
R12685 VSS.n4130 VSS.n4129 9.3
R12686 VSS.n4342 VSS.n4341 9.3
R12687 VSS.n4341 VSS.n4340 9.3
R12688 VSS.n4340 VSS.n4339 9.3
R12689 VSS.n4343 VSS.n4117 9.3
R12690 VSS.n4346 VSS.n4112 9.3
R12691 VSS.n4347 VSS.n4346 9.3
R12692 VSS.n4348 VSS.n4347 9.3
R12693 VSS.n4354 VSS.n4353 9.3
R12694 VSS.n4357 VSS.n4356 9.3
R12695 VSS.n4357 VSS.n4107 9.3
R12696 VSS.n4107 VSS.n4106 9.3
R12697 VSS.n4111 VSS.n4110 9.3
R12698 VSS.n4365 VSS.n4364 9.3
R12699 VSS.n4364 VSS.n4363 9.3
R12700 VSS.n4363 VSS.n4362 9.3
R12701 VSS.n4366 VSS.n4098 9.3
R12702 VSS.n4369 VSS.n4093 9.3
R12703 VSS.n4370 VSS.n4369 9.3
R12704 VSS.n4371 VSS.n4370 9.3
R12705 VSS.n4377 VSS.n4376 9.3
R12706 VSS.n4380 VSS.n4379 9.3
R12707 VSS.n4380 VSS.n4088 9.3
R12708 VSS.n4088 VSS.n4087 9.3
R12709 VSS.n4092 VSS.n4091 9.3
R12710 VSS.n4388 VSS.n4387 9.3
R12711 VSS.n4387 VSS.n4386 9.3
R12712 VSS.n4386 VSS.n4385 9.3
R12713 VSS.n4389 VSS.n4079 9.3
R12714 VSS.n4392 VSS.n4074 9.3
R12715 VSS.n4393 VSS.n4392 9.3
R12716 VSS.n4394 VSS.n4393 9.3
R12717 VSS.n4400 VSS.n4399 9.3
R12718 VSS.n4403 VSS.n4402 9.3
R12719 VSS.n4403 VSS.n4069 9.3
R12720 VSS.n4069 VSS.n4068 9.3
R12721 VSS.n4073 VSS.n4072 9.3
R12722 VSS.n4411 VSS.n4410 9.3
R12723 VSS.n4410 VSS.n4409 9.3
R12724 VSS.n4409 VSS.n4408 9.3
R12725 VSS.n4414 VSS.n4413 9.3
R12726 VSS.n4417 VSS.n4416 9.3
R12727 VSS.n4418 VSS.n4417 9.3
R12728 VSS.n4419 VSS.n4418 9.3
R12729 VSS.n4059 VSS.n4058 9.3
R12730 VSS.n4050 VSS.n4049 9.3
R12731 VSS.n4050 VSS.n3329 9.3
R12732 VSS.n4054 VSS.n3329 9.3
R12733 VSS.n4048 VSS.n4047 9.3
R12734 VSS.n4045 VSS.n3335 9.3
R12735 VSS.n4045 VSS.n4044 9.3
R12736 VSS.n4044 VSS.n4043 9.3
R12737 VSS.n4038 VSS.n4037 9.3
R12738 VSS.n4035 VSS.n4034 9.3
R12739 VSS.n4034 VSS.n3338 9.3
R12740 VSS.n3338 VSS.n3337 9.3
R12741 VSS.n3346 VSS.n3340 9.3
R12742 VSS.n4027 VSS.n4026 9.3
R12743 VSS.n4028 VSS.n4027 9.3
R12744 VSS.n4029 VSS.n4028 9.3
R12745 VSS.n4024 VSS.n4023 9.3
R12746 VSS.n4015 VSS.n4014 9.3
R12747 VSS.n4015 VSS.n3350 9.3
R12748 VSS.n4019 VSS.n3350 9.3
R12749 VSS.n4013 VSS.n4012 9.3
R12750 VSS.n4010 VSS.n3356 9.3
R12751 VSS.n4010 VSS.n4009 9.3
R12752 VSS.n4009 VSS.n4008 9.3
R12753 VSS.n4003 VSS.n4002 9.3
R12754 VSS.n4000 VSS.n3999 9.3
R12755 VSS.n3999 VSS.n3359 9.3
R12756 VSS.n3359 VSS.n3358 9.3
R12757 VSS.n3367 VSS.n3361 9.3
R12758 VSS.n3992 VSS.n3991 9.3
R12759 VSS.n3993 VSS.n3992 9.3
R12760 VSS.n3994 VSS.n3993 9.3
R12761 VSS.n3989 VSS.n3988 9.3
R12762 VSS.n3980 VSS.n3979 9.3
R12763 VSS.n3980 VSS.n3371 9.3
R12764 VSS.n3984 VSS.n3371 9.3
R12765 VSS.n3978 VSS.n3977 9.3
R12766 VSS.n3975 VSS.n3377 9.3
R12767 VSS.n3975 VSS.n3974 9.3
R12768 VSS.n3974 VSS.n3973 9.3
R12769 VSS.n3968 VSS.n3967 9.3
R12770 VSS.n3965 VSS.n3964 9.3
R12771 VSS.n3964 VSS.n3380 9.3
R12772 VSS.n3380 VSS.n3379 9.3
R12773 VSS.n3953 VSS.n3952 9.3
R12774 VSS.n3956 VSS.n3955 9.3
R12775 VSS.n3957 VSS.n3956 9.3
R12776 VSS.n3958 VSS.n3957 9.3
R12777 VSS.n3631 VSS.n3391 9.3
R12778 VSS.n3637 VSS.n3636 9.3
R12779 VSS.n3637 VSS.n3626 9.3
R12780 VSS.n3626 VSS.n3625 9.3
R12781 VSS.n3634 VSS.n3633 9.3
R12782 VSS.n3645 VSS.n3644 9.3
R12783 VSS.n3644 VSS.n3643 9.3
R12784 VSS.n3643 VSS.n3642 9.3
R12785 VSS.n3646 VSS.n3617 9.3
R12786 VSS.n3649 VSS.n3612 9.3
R12787 VSS.n3650 VSS.n3649 9.3
R12788 VSS.n3651 VSS.n3650 9.3
R12789 VSS.n3657 VSS.n3656 9.3
R12790 VSS.n3660 VSS.n3659 9.3
R12791 VSS.n3660 VSS.n3607 9.3
R12792 VSS.n3607 VSS.n3606 9.3
R12793 VSS.n3611 VSS.n3610 9.3
R12794 VSS.n3668 VSS.n3667 9.3
R12795 VSS.n3667 VSS.n3666 9.3
R12796 VSS.n3666 VSS.n3665 9.3
R12797 VSS.n3669 VSS.n3598 9.3
R12798 VSS.n3672 VSS.n3593 9.3
R12799 VSS.n3673 VSS.n3672 9.3
R12800 VSS.n3674 VSS.n3673 9.3
R12801 VSS.n3680 VSS.n3679 9.3
R12802 VSS.n3683 VSS.n3682 9.3
R12803 VSS.n3683 VSS.n3588 9.3
R12804 VSS.n3588 VSS.n3587 9.3
R12805 VSS.n3592 VSS.n3591 9.3
R12806 VSS.n3691 VSS.n3690 9.3
R12807 VSS.n3690 VSS.n3689 9.3
R12808 VSS.n3689 VSS.n3688 9.3
R12809 VSS.n3692 VSS.n3579 9.3
R12810 VSS.n3695 VSS.n3574 9.3
R12811 VSS.n3696 VSS.n3695 9.3
R12812 VSS.n3697 VSS.n3696 9.3
R12813 VSS.n3703 VSS.n3702 9.3
R12814 VSS.n3706 VSS.n3705 9.3
R12815 VSS.n3706 VSS.n3569 9.3
R12816 VSS.n3569 VSS.n3568 9.3
R12817 VSS.n3573 VSS.n3572 9.3
R12818 VSS.n3714 VSS.n3713 9.3
R12819 VSS.n3713 VSS.n3712 9.3
R12820 VSS.n3712 VSS.n3711 9.3
R12821 VSS.n3716 VSS.n3524 9.3
R12822 VSS.n3719 VSS.n3519 9.3
R12823 VSS.n3720 VSS.n3719 9.3
R12824 VSS.n3721 VSS.n3720 9.3
R12825 VSS.n3727 VSS.n3726 9.3
R12826 VSS.n3730 VSS.n3729 9.3
R12827 VSS.n3730 VSS.n3514 9.3
R12828 VSS.n3514 VSS.n3513 9.3
R12829 VSS.n3518 VSS.n3517 9.3
R12830 VSS.n3738 VSS.n3737 9.3
R12831 VSS.n3737 VSS.n3736 9.3
R12832 VSS.n3736 VSS.n3735 9.3
R12833 VSS.n3739 VSS.n3505 9.3
R12834 VSS.n3742 VSS.n3500 9.3
R12835 VSS.n3743 VSS.n3742 9.3
R12836 VSS.n3744 VSS.n3743 9.3
R12837 VSS.n3750 VSS.n3749 9.3
R12838 VSS.n3753 VSS.n3752 9.3
R12839 VSS.n3753 VSS.n3495 9.3
R12840 VSS.n3495 VSS.n3494 9.3
R12841 VSS.n3499 VSS.n3498 9.3
R12842 VSS.n3761 VSS.n3760 9.3
R12843 VSS.n3760 VSS.n3759 9.3
R12844 VSS.n3759 VSS.n3758 9.3
R12845 VSS.n3762 VSS.n3486 9.3
R12846 VSS.n3765 VSS.n3481 9.3
R12847 VSS.n3766 VSS.n3765 9.3
R12848 VSS.n3767 VSS.n3766 9.3
R12849 VSS.n3773 VSS.n3772 9.3
R12850 VSS.n3776 VSS.n3775 9.3
R12851 VSS.n3776 VSS.n3476 9.3
R12852 VSS.n3476 VSS.n3475 9.3
R12853 VSS.n3480 VSS.n3479 9.3
R12854 VSS.n3784 VSS.n3783 9.3
R12855 VSS.n3783 VSS.n3782 9.3
R12856 VSS.n3782 VSS.n3781 9.3
R12857 VSS.n3785 VSS.n3467 9.3
R12858 VSS.n3788 VSS.n3462 9.3
R12859 VSS.n3789 VSS.n3788 9.3
R12860 VSS.n3790 VSS.n3789 9.3
R12861 VSS.n3796 VSS.n3795 9.3
R12862 VSS.n3799 VSS.n3798 9.3
R12863 VSS.n3799 VSS.n3456 9.3
R12864 VSS.n3456 VSS.n3455 9.3
R12865 VSS.n3461 VSS.n3460 9.3
R12866 VSS.n3806 VSS.n3453 9.3
R12867 VSS.n3806 VSS.n3805 9.3
R12868 VSS.n3805 VSS.n3804 9.3
R12869 VSS.n4839 VSS.n4833 9.3
R12870 VSS.n4840 VSS.n4839 9.3
R12871 VSS.n4841 VSS.n4840 9.3
R12872 VSS.n4836 VSS.n3095 9.3
R12873 VSS.n3040 VSS.n3039 9.3
R12874 VSS.n3039 VSS.n1658 9.3
R12875 VSS.n3088 VSS.n1658 9.3
R12876 VSS.n3051 VSS.n3050 9.3
R12877 VSS.n3050 VSS.n1683 9.3
R12878 VSS.n3053 VSS.n3052 9.3
R12879 VSS.n3057 VSS.n3056 9.3
R12880 VSS.n3056 VSS.n3055 9.3
R12881 VSS.n3063 VSS.n3062 9.3
R12882 VSS.n3062 VSS.n3061 9.3
R12883 VSS.n3065 VSS.n3064 9.3
R12884 VSS.n3069 VSS.n3068 9.3
R12885 VSS.n3068 VSS.n3067 9.3
R12886 VSS.n3074 VSS.n3013 9.3
R12887 VSS.n3074 VSS.n3073 9.3
R12888 VSS.n3079 VSS.n3078 9.3
R12889 VSS.n3083 VSS.n3081 9.3
R12890 VSS.n3083 VSS.n3082 9.3
R12891 VSS.n3009 VSS.n1696 9.3
R12892 VSS.n3009 VSS.n1693 9.3
R12893 VSS.n3012 VSS.n1694 9.3
R12894 VSS.n3048 VSS.n3047 9.3
R12895 VSS.n3059 VSS.n3058 9.3
R12896 VSS.n3070 VSS.n3014 9.3
R12897 VSS.n2950 VSS.n2949 9.3
R12898 VSS.n2949 VSS.n1748 9.3
R12899 VSS.n2998 VSS.n1748 9.3
R12900 VSS.n2961 VSS.n2960 9.3
R12901 VSS.n2960 VSS.n1773 9.3
R12902 VSS.n2963 VSS.n2962 9.3
R12903 VSS.n2967 VSS.n2966 9.3
R12904 VSS.n2966 VSS.n2965 9.3
R12905 VSS.n2973 VSS.n2972 9.3
R12906 VSS.n2972 VSS.n2971 9.3
R12907 VSS.n2975 VSS.n2974 9.3
R12908 VSS.n2979 VSS.n2978 9.3
R12909 VSS.n2978 VSS.n2977 9.3
R12910 VSS.n2984 VSS.n2923 9.3
R12911 VSS.n2984 VSS.n2983 9.3
R12912 VSS.n2989 VSS.n2988 9.3
R12913 VSS.n2993 VSS.n2991 9.3
R12914 VSS.n2993 VSS.n2992 9.3
R12915 VSS.n2919 VSS.n1786 9.3
R12916 VSS.n2919 VSS.n1783 9.3
R12917 VSS.n2922 VSS.n1784 9.3
R12918 VSS.n2958 VSS.n2957 9.3
R12919 VSS.n2969 VSS.n2968 9.3
R12920 VSS.n2980 VSS.n2924 9.3
R12921 VSS.n2860 VSS.n2859 9.3
R12922 VSS.n2859 VSS.n1838 9.3
R12923 VSS.n2908 VSS.n1838 9.3
R12924 VSS.n2871 VSS.n2870 9.3
R12925 VSS.n2870 VSS.n1863 9.3
R12926 VSS.n2873 VSS.n2872 9.3
R12927 VSS.n2877 VSS.n2876 9.3
R12928 VSS.n2876 VSS.n2875 9.3
R12929 VSS.n2883 VSS.n2882 9.3
R12930 VSS.n2882 VSS.n2881 9.3
R12931 VSS.n2885 VSS.n2884 9.3
R12932 VSS.n2889 VSS.n2888 9.3
R12933 VSS.n2888 VSS.n2887 9.3
R12934 VSS.n2894 VSS.n2833 9.3
R12935 VSS.n2894 VSS.n2893 9.3
R12936 VSS.n2899 VSS.n2898 9.3
R12937 VSS.n2903 VSS.n2901 9.3
R12938 VSS.n2903 VSS.n2902 9.3
R12939 VSS.n2829 VSS.n1876 9.3
R12940 VSS.n2829 VSS.n1873 9.3
R12941 VSS.n2832 VSS.n1874 9.3
R12942 VSS.n2868 VSS.n2867 9.3
R12943 VSS.n2879 VSS.n2878 9.3
R12944 VSS.n2890 VSS.n2834 9.3
R12945 VSS.n2770 VSS.n2769 9.3
R12946 VSS.n2769 VSS.n1928 9.3
R12947 VSS.n2818 VSS.n1928 9.3
R12948 VSS.n2781 VSS.n2780 9.3
R12949 VSS.n2780 VSS.n1953 9.3
R12950 VSS.n2783 VSS.n2782 9.3
R12951 VSS.n2787 VSS.n2786 9.3
R12952 VSS.n2786 VSS.n2785 9.3
R12953 VSS.n2793 VSS.n2792 9.3
R12954 VSS.n2792 VSS.n2791 9.3
R12955 VSS.n2795 VSS.n2794 9.3
R12956 VSS.n2799 VSS.n2798 9.3
R12957 VSS.n2798 VSS.n2797 9.3
R12958 VSS.n2804 VSS.n2743 9.3
R12959 VSS.n2804 VSS.n2803 9.3
R12960 VSS.n2809 VSS.n2808 9.3
R12961 VSS.n2813 VSS.n2811 9.3
R12962 VSS.n2813 VSS.n2812 9.3
R12963 VSS.n2739 VSS.n1966 9.3
R12964 VSS.n2739 VSS.n1963 9.3
R12965 VSS.n2742 VSS.n1964 9.3
R12966 VSS.n2778 VSS.n2777 9.3
R12967 VSS.n2789 VSS.n2788 9.3
R12968 VSS.n2800 VSS.n2744 9.3
R12969 VSS.n2680 VSS.n2679 9.3
R12970 VSS.n2679 VSS.n2018 9.3
R12971 VSS.n2728 VSS.n2018 9.3
R12972 VSS.n2691 VSS.n2690 9.3
R12973 VSS.n2690 VSS.n2043 9.3
R12974 VSS.n2693 VSS.n2692 9.3
R12975 VSS.n2697 VSS.n2696 9.3
R12976 VSS.n2696 VSS.n2695 9.3
R12977 VSS.n2703 VSS.n2702 9.3
R12978 VSS.n2702 VSS.n2701 9.3
R12979 VSS.n2705 VSS.n2704 9.3
R12980 VSS.n2709 VSS.n2708 9.3
R12981 VSS.n2708 VSS.n2707 9.3
R12982 VSS.n2714 VSS.n2653 9.3
R12983 VSS.n2714 VSS.n2713 9.3
R12984 VSS.n2719 VSS.n2718 9.3
R12985 VSS.n2723 VSS.n2721 9.3
R12986 VSS.n2723 VSS.n2722 9.3
R12987 VSS.n2649 VSS.n2056 9.3
R12988 VSS.n2649 VSS.n2053 9.3
R12989 VSS.n2652 VSS.n2054 9.3
R12990 VSS.n2688 VSS.n2687 9.3
R12991 VSS.n2699 VSS.n2698 9.3
R12992 VSS.n2710 VSS.n2654 9.3
R12993 VSS.n2590 VSS.n2589 9.3
R12994 VSS.n2589 VSS.n2108 9.3
R12995 VSS.n2638 VSS.n2108 9.3
R12996 VSS.n2601 VSS.n2600 9.3
R12997 VSS.n2600 VSS.n2133 9.3
R12998 VSS.n2603 VSS.n2602 9.3
R12999 VSS.n2607 VSS.n2606 9.3
R13000 VSS.n2606 VSS.n2605 9.3
R13001 VSS.n2613 VSS.n2612 9.3
R13002 VSS.n2612 VSS.n2611 9.3
R13003 VSS.n2615 VSS.n2614 9.3
R13004 VSS.n2619 VSS.n2618 9.3
R13005 VSS.n2618 VSS.n2617 9.3
R13006 VSS.n2624 VSS.n2563 9.3
R13007 VSS.n2624 VSS.n2623 9.3
R13008 VSS.n2629 VSS.n2628 9.3
R13009 VSS.n2633 VSS.n2631 9.3
R13010 VSS.n2633 VSS.n2632 9.3
R13011 VSS.n2559 VSS.n2146 9.3
R13012 VSS.n2559 VSS.n2143 9.3
R13013 VSS.n2562 VSS.n2144 9.3
R13014 VSS.n2598 VSS.n2597 9.3
R13015 VSS.n2609 VSS.n2608 9.3
R13016 VSS.n2620 VSS.n2564 9.3
R13017 VSS.n2500 VSS.n2499 9.3
R13018 VSS.n2499 VSS.n2198 9.3
R13019 VSS.n2548 VSS.n2198 9.3
R13020 VSS.n2511 VSS.n2510 9.3
R13021 VSS.n2510 VSS.n2223 9.3
R13022 VSS.n2513 VSS.n2512 9.3
R13023 VSS.n2517 VSS.n2516 9.3
R13024 VSS.n2516 VSS.n2515 9.3
R13025 VSS.n2523 VSS.n2522 9.3
R13026 VSS.n2522 VSS.n2521 9.3
R13027 VSS.n2525 VSS.n2524 9.3
R13028 VSS.n2529 VSS.n2528 9.3
R13029 VSS.n2528 VSS.n2527 9.3
R13030 VSS.n2534 VSS.n2473 9.3
R13031 VSS.n2534 VSS.n2533 9.3
R13032 VSS.n2539 VSS.n2538 9.3
R13033 VSS.n2543 VSS.n2541 9.3
R13034 VSS.n2543 VSS.n2542 9.3
R13035 VSS.n2469 VSS.n2236 9.3
R13036 VSS.n2469 VSS.n2233 9.3
R13037 VSS.n2472 VSS.n2234 9.3
R13038 VSS.n2508 VSS.n2507 9.3
R13039 VSS.n2519 VSS.n2518 9.3
R13040 VSS.n2530 VSS.n2474 9.3
R13041 VSS.n2410 VSS.n2409 9.3
R13042 VSS.n2409 VSS.n2288 9.3
R13043 VSS.n2458 VSS.n2288 9.3
R13044 VSS.n2421 VSS.n2420 9.3
R13045 VSS.n2420 VSS.n2313 9.3
R13046 VSS.n2423 VSS.n2422 9.3
R13047 VSS.n2427 VSS.n2426 9.3
R13048 VSS.n2426 VSS.n2425 9.3
R13049 VSS.n2433 VSS.n2432 9.3
R13050 VSS.n2432 VSS.n2431 9.3
R13051 VSS.n2435 VSS.n2434 9.3
R13052 VSS.n2439 VSS.n2438 9.3
R13053 VSS.n2438 VSS.n2437 9.3
R13054 VSS.n2444 VSS.n2383 9.3
R13055 VSS.n2444 VSS.n2443 9.3
R13056 VSS.n2449 VSS.n2448 9.3
R13057 VSS.n2453 VSS.n2451 9.3
R13058 VSS.n2453 VSS.n2452 9.3
R13059 VSS.n2379 VSS.n2326 9.3
R13060 VSS.n2379 VSS.n2323 9.3
R13061 VSS.n2382 VSS.n2324 9.3
R13062 VSS.n2418 VSS.n2417 9.3
R13063 VSS.n2429 VSS.n2428 9.3
R13064 VSS.n2440 VSS.n2384 9.3
R13065 VSS.n2416 VSS.n2415 9.3
R13066 VSS.n2415 VSS.n2414 9.3
R13067 VSS.n2412 VSS.n2411 9.3
R13068 VSS.n2286 VSS.n2285 9.3
R13069 VSS.n2506 VSS.n2505 9.3
R13070 VSS.n2505 VSS.n2504 9.3
R13071 VSS.n2502 VSS.n2501 9.3
R13072 VSS.n2196 VSS.n2195 9.3
R13073 VSS.n2596 VSS.n2595 9.3
R13074 VSS.n2595 VSS.n2594 9.3
R13075 VSS.n2592 VSS.n2591 9.3
R13076 VSS.n2106 VSS.n2105 9.3
R13077 VSS.n2686 VSS.n2685 9.3
R13078 VSS.n2685 VSS.n2684 9.3
R13079 VSS.n2682 VSS.n2681 9.3
R13080 VSS.n2016 VSS.n2015 9.3
R13081 VSS.n2776 VSS.n2775 9.3
R13082 VSS.n2775 VSS.n2774 9.3
R13083 VSS.n2772 VSS.n2771 9.3
R13084 VSS.n1926 VSS.n1925 9.3
R13085 VSS.n2866 VSS.n2865 9.3
R13086 VSS.n2865 VSS.n2864 9.3
R13087 VSS.n2862 VSS.n2861 9.3
R13088 VSS.n1836 VSS.n1835 9.3
R13089 VSS.n2956 VSS.n2955 9.3
R13090 VSS.n2955 VSS.n2954 9.3
R13091 VSS.n2952 VSS.n2951 9.3
R13092 VSS.n1746 VSS.n1745 9.3
R13093 VSS.n3046 VSS.n3045 9.3
R13094 VSS.n3045 VSS.n3044 9.3
R13095 VSS.n3042 VSS.n3041 9.3
R13096 VSS.n1656 VSS.n1655 9.3
R13097 VSS.n1183 VSS.n1182 9.3
R13098 VSS.n1183 VSS.n1084 9.3
R13099 VSS.n1084 VSS.n1083 9.3
R13100 VSS.n1088 VSS.n1087 9.3
R13101 VSS.n1191 VSS.n1190 9.3
R13102 VSS.n1190 VSS.n1189 9.3
R13103 VSS.n1189 VSS.n1188 9.3
R13104 VSS.n1195 VSS.n1070 9.3
R13105 VSS.n1196 VSS.n1195 9.3
R13106 VSS.n1197 VSS.n1196 9.3
R13107 VSS.n1203 VSS.n1202 9.3
R13108 VSS.n1206 VSS.n1205 9.3
R13109 VSS.n1206 VSS.n1065 9.3
R13110 VSS.n1065 VSS.n1064 9.3
R13111 VSS.n1214 VSS.n1213 9.3
R13112 VSS.n1213 VSS.n1212 9.3
R13113 VSS.n1212 VSS.n1211 9.3
R13114 VSS.n1215 VSS.n1056 9.3
R13115 VSS.n1218 VSS.n1051 9.3
R13116 VSS.n1219 VSS.n1218 9.3
R13117 VSS.n1220 VSS.n1219 9.3
R13118 VSS.n1229 VSS.n1228 9.3
R13119 VSS.n1229 VSS.n1046 9.3
R13120 VSS.n1046 VSS.n1045 9.3
R13121 VSS.n1050 VSS.n1049 9.3
R13122 VSS.n1237 VSS.n1236 9.3
R13123 VSS.n1236 VSS.n1235 9.3
R13124 VSS.n1235 VSS.n1234 9.3
R13125 VSS.n1241 VSS.n1032 9.3
R13126 VSS.n1242 VSS.n1241 9.3
R13127 VSS.n1243 VSS.n1242 9.3
R13128 VSS.n1249 VSS.n1248 9.3
R13129 VSS.n1252 VSS.n1251 9.3
R13130 VSS.n1252 VSS.n1027 9.3
R13131 VSS.n1027 VSS.n1026 9.3
R13132 VSS.n1260 VSS.n1259 9.3
R13133 VSS.n1259 VSS.n1258 9.3
R13134 VSS.n1258 VSS.n1257 9.3
R13135 VSS.n1180 VSS.n1179 9.3
R13136 VSS.n1192 VSS.n1075 9.3
R13137 VSS.n1069 VSS.n1068 9.3
R13138 VSS.n1226 VSS.n1225 9.3
R13139 VSS.n1238 VSS.n1037 9.3
R13140 VSS.n1031 VSS.n1030 9.3
R13141 VSS.n1263 VSS.n1262 9.3
R13142 VSS.n1266 VSS.n1265 9.3
R13143 VSS.n1267 VSS.n1266 9.3
R13144 VSS.n1268 VSS.n1267 9.3
R13145 VSS.n1017 VSS.n1016 9.3
R13146 VSS.n1008 VSS.n1007 9.3
R13147 VSS.n1008 VSS.n659 9.3
R13148 VSS.n1012 VSS.n659 9.3
R13149 VSS.n1006 VSS.n1005 9.3
R13150 VSS.n1003 VSS.n665 9.3
R13151 VSS.n1003 VSS.n1002 9.3
R13152 VSS.n1002 VSS.n1001 9.3
R13153 VSS.n996 VSS.n995 9.3
R13154 VSS.n993 VSS.n992 9.3
R13155 VSS.n992 VSS.n668 9.3
R13156 VSS.n668 VSS.n667 9.3
R13157 VSS.n676 VSS.n670 9.3
R13158 VSS.n985 VSS.n984 9.3
R13159 VSS.n986 VSS.n985 9.3
R13160 VSS.n987 VSS.n986 9.3
R13161 VSS.n982 VSS.n981 9.3
R13162 VSS.n973 VSS.n972 9.3
R13163 VSS.n973 VSS.n680 9.3
R13164 VSS.n977 VSS.n680 9.3
R13165 VSS.n971 VSS.n970 9.3
R13166 VSS.n968 VSS.n686 9.3
R13167 VSS.n968 VSS.n967 9.3
R13168 VSS.n967 VSS.n966 9.3
R13169 VSS.n961 VSS.n960 9.3
R13170 VSS.n958 VSS.n957 9.3
R13171 VSS.n957 VSS.n689 9.3
R13172 VSS.n689 VSS.n688 9.3
R13173 VSS.n697 VSS.n691 9.3
R13174 VSS.n950 VSS.n949 9.3
R13175 VSS.n951 VSS.n950 9.3
R13176 VSS.n952 VSS.n951 9.3
R13177 VSS.n947 VSS.n946 9.3
R13178 VSS.n938 VSS.n937 9.3
R13179 VSS.n938 VSS.n701 9.3
R13180 VSS.n942 VSS.n701 9.3
R13181 VSS.n936 VSS.n935 9.3
R13182 VSS.n933 VSS.n707 9.3
R13183 VSS.n933 VSS.n932 9.3
R13184 VSS.n932 VSS.n931 9.3
R13185 VSS.n926 VSS.n925 9.3
R13186 VSS.n923 VSS.n922 9.3
R13187 VSS.n922 VSS.n710 9.3
R13188 VSS.n710 VSS.n709 9.3
R13189 VSS.n884 VSS.n883 9.3
R13190 VSS.n881 VSS.n880 9.3
R13191 VSS.n880 VSS.n879 9.3
R13192 VSS.n879 VSS.n715 9.3
R13193 VSS.n727 VSS.n720 9.3
R13194 VSS.n873 VSS.n872 9.3
R13195 VSS.n874 VSS.n873 9.3
R13196 VSS.n875 VSS.n874 9.3
R13197 VSS.n870 VSS.n869 9.3
R13198 VSS.n861 VSS.n860 9.3
R13199 VSS.n861 VSS.n731 9.3
R13200 VSS.n865 VSS.n731 9.3
R13201 VSS.n859 VSS.n858 9.3
R13202 VSS.n856 VSS.n737 9.3
R13203 VSS.n856 VSS.n855 9.3
R13204 VSS.n855 VSS.n854 9.3
R13205 VSS.n849 VSS.n848 9.3
R13206 VSS.n846 VSS.n845 9.3
R13207 VSS.n845 VSS.n740 9.3
R13208 VSS.n740 VSS.n739 9.3
R13209 VSS.n748 VSS.n742 9.3
R13210 VSS.n838 VSS.n837 9.3
R13211 VSS.n839 VSS.n838 9.3
R13212 VSS.n840 VSS.n839 9.3
R13213 VSS.n835 VSS.n834 9.3
R13214 VSS.n826 VSS.n825 9.3
R13215 VSS.n826 VSS.n752 9.3
R13216 VSS.n830 VSS.n752 9.3
R13217 VSS.n824 VSS.n823 9.3
R13218 VSS.n821 VSS.n758 9.3
R13219 VSS.n821 VSS.n820 9.3
R13220 VSS.n820 VSS.n819 9.3
R13221 VSS.n814 VSS.n813 9.3
R13222 VSS.n811 VSS.n810 9.3
R13223 VSS.n810 VSS.n761 9.3
R13224 VSS.n761 VSS.n760 9.3
R13225 VSS.n769 VSS.n763 9.3
R13226 VSS.n803 VSS.n802 9.3
R13227 VSS.n804 VSS.n803 9.3
R13228 VSS.n805 VSS.n804 9.3
R13229 VSS.n800 VSS.n799 9.3
R13230 VSS.n791 VSS.n790 9.3
R13231 VSS.n791 VSS.n773 9.3
R13232 VSS.n795 VSS.n773 9.3
R13233 VSS.n789 VSS.n788 9.3
R13234 VSS.n786 VSS.n779 9.3
R13235 VSS.n786 VSS.n785 9.3
R13236 VSS.n785 VSS.n784 9.3
R13237 VSS.n5703 VSS.n5702 9.3
R13238 VSS.n5706 VSS.n5705 9.3
R13239 VSS.n5706 VSS.n584 9.3
R13240 VSS.n584 VSS.n583 9.3
R13241 VSS.n588 VSS.n587 9.3
R13242 VSS.n5714 VSS.n5713 9.3
R13243 VSS.n5713 VSS.n5712 9.3
R13244 VSS.n5712 VSS.n5711 9.3
R13245 VSS.n5715 VSS.n575 9.3
R13246 VSS.n5718 VSS.n570 9.3
R13247 VSS.n5719 VSS.n5718 9.3
R13248 VSS.n5720 VSS.n5719 9.3
R13249 VSS.n5726 VSS.n5725 9.3
R13250 VSS.n5729 VSS.n5728 9.3
R13251 VSS.n5729 VSS.n565 9.3
R13252 VSS.n565 VSS.n564 9.3
R13253 VSS.n569 VSS.n568 9.3
R13254 VSS.n5737 VSS.n5736 9.3
R13255 VSS.n5736 VSS.n5735 9.3
R13256 VSS.n5735 VSS.n5734 9.3
R13257 VSS.n5738 VSS.n556 9.3
R13258 VSS.n5741 VSS.n551 9.3
R13259 VSS.n5742 VSS.n5741 9.3
R13260 VSS.n5743 VSS.n5742 9.3
R13261 VSS.n5749 VSS.n5748 9.3
R13262 VSS.n5752 VSS.n5751 9.3
R13263 VSS.n5752 VSS.n546 9.3
R13264 VSS.n546 VSS.n545 9.3
R13265 VSS.n550 VSS.n549 9.3
R13266 VSS.n5760 VSS.n5759 9.3
R13267 VSS.n5759 VSS.n5758 9.3
R13268 VSS.n5758 VSS.n5757 9.3
R13269 VSS.n5761 VSS.n537 9.3
R13270 VSS.n5764 VSS.n532 9.3
R13271 VSS.n5765 VSS.n5764 9.3
R13272 VSS.n5766 VSS.n5765 9.3
R13273 VSS.n5772 VSS.n5771 9.3
R13274 VSS.n5775 VSS.n5774 9.3
R13275 VSS.n5775 VSS.n527 9.3
R13276 VSS.n527 VSS.n526 9.3
R13277 VSS.n531 VSS.n530 9.3
R13278 VSS.n5783 VSS.n5782 9.3
R13279 VSS.n5782 VSS.n5781 9.3
R13280 VSS.n5781 VSS.n5780 9.3
R13281 VSS.n5600 VSS.n519 9.3
R13282 VSS.n5604 VSS.n5603 9.3
R13283 VSS.n5604 VSS.n5595 9.3
R13284 VSS.n5596 VSS.n5595 9.3
R13285 VSS.n5616 VSS.n5615 9.3
R13286 VSS.n5613 VSS.n5612 9.3
R13287 VSS.n5612 VSS.n5611 9.3
R13288 VSS.n5611 VSS.n5610 9.3
R13289 VSS.n5589 VSS.n1383 9.3
R13290 VSS.n5586 VSS.n1389 9.3
R13291 VSS.n1389 VSS.n1388 9.3
R13292 VSS.n1388 VSS.n1387 9.3
R13293 VSS.n5585 VSS.n5584 9.3
R13294 VSS.n5575 VSS.n5574 9.3
R13295 VSS.n5575 VSS.n1393 9.3
R13296 VSS.n5579 VSS.n1393 9.3
R13297 VSS.n5573 VSS.n5572 9.3
R13298 VSS.n5570 VSS.n1400 9.3
R13299 VSS.n5570 VSS.n5569 9.3
R13300 VSS.n5569 VSS.n5568 9.3
R13301 VSS.n5563 VSS.n5562 9.3
R13302 VSS.n5560 VSS.n5559 9.3
R13303 VSS.n5559 VSS.n1403 9.3
R13304 VSS.n1403 VSS.n1402 9.3
R13305 VSS.n1411 VSS.n1405 9.3
R13306 VSS.n5552 VSS.n5551 9.3
R13307 VSS.n5553 VSS.n5552 9.3
R13308 VSS.n5554 VSS.n5553 9.3
R13309 VSS.n5549 VSS.n5548 9.3
R13310 VSS.n5540 VSS.n5539 9.3
R13311 VSS.n5540 VSS.n1415 9.3
R13312 VSS.n5544 VSS.n1415 9.3
R13313 VSS.n5538 VSS.n5537 9.3
R13314 VSS.n5535 VSS.n1421 9.3
R13315 VSS.n5535 VSS.n5534 9.3
R13316 VSS.n5534 VSS.n5533 9.3
R13317 VSS.n5528 VSS.n5527 9.3
R13318 VSS.n5525 VSS.n5524 9.3
R13319 VSS.n5524 VSS.n1424 9.3
R13320 VSS.n1424 VSS.n1423 9.3
R13321 VSS.n1432 VSS.n1426 9.3
R13322 VSS.n5517 VSS.n5516 9.3
R13323 VSS.n5518 VSS.n5517 9.3
R13324 VSS.n5519 VSS.n5518 9.3
R13325 VSS.n5514 VSS.n5513 9.3
R13326 VSS.n5505 VSS.n5504 9.3
R13327 VSS.n5505 VSS.n1436 9.3
R13328 VSS.n5509 VSS.n1436 9.3
R13329 VSS.n5503 VSS.n5502 9.3
R13330 VSS.n5500 VSS.n1442 9.3
R13331 VSS.n5500 VSS.n5499 9.3
R13332 VSS.n5499 VSS.n5498 9.3
R13333 VSS.n5302 VSS.n1446 9.3
R13334 VSS.n5312 VSS.n5311 9.3
R13335 VSS.n5311 VSS.n5310 9.3
R13336 VSS.n5310 VSS.n5309 9.3
R13337 VSS.n5313 VSS.n5301 9.3
R13338 VSS.n5316 VSS.n5296 9.3
R13339 VSS.n5317 VSS.n5316 9.3
R13340 VSS.n5318 VSS.n5317 9.3
R13341 VSS.n5324 VSS.n5323 9.3
R13342 VSS.n5327 VSS.n5326 9.3
R13343 VSS.n5327 VSS.n5291 9.3
R13344 VSS.n5291 VSS.n5290 9.3
R13345 VSS.n5295 VSS.n5294 9.3
R13346 VSS.n5335 VSS.n5334 9.3
R13347 VSS.n5334 VSS.n5333 9.3
R13348 VSS.n5333 VSS.n5332 9.3
R13349 VSS.n5336 VSS.n5282 9.3
R13350 VSS.n5339 VSS.n5277 9.3
R13351 VSS.n5340 VSS.n5339 9.3
R13352 VSS.n5341 VSS.n5340 9.3
R13353 VSS.n5347 VSS.n5346 9.3
R13354 VSS.n5350 VSS.n5349 9.3
R13355 VSS.n5350 VSS.n5272 9.3
R13356 VSS.n5272 VSS.n5271 9.3
R13357 VSS.n5276 VSS.n5275 9.3
R13358 VSS.n5358 VSS.n5357 9.3
R13359 VSS.n5357 VSS.n5356 9.3
R13360 VSS.n5356 VSS.n5355 9.3
R13361 VSS.n5359 VSS.n5263 9.3
R13362 VSS.n5362 VSS.n5258 9.3
R13363 VSS.n5363 VSS.n5362 9.3
R13364 VSS.n5364 VSS.n5363 9.3
R13365 VSS.n5370 VSS.n5369 9.3
R13366 VSS.n5373 VSS.n5372 9.3
R13367 VSS.n5373 VSS.n5253 9.3
R13368 VSS.n5253 VSS.n5252 9.3
R13369 VSS.n5257 VSS.n5256 9.3
R13370 VSS.n5381 VSS.n5380 9.3
R13371 VSS.n5380 VSS.n5379 9.3
R13372 VSS.n5379 VSS.n5378 9.3
R13373 VSS.n5382 VSS.n5244 9.3
R13374 VSS.n5385 VSS.n5238 9.3
R13375 VSS.n5386 VSS.n5385 9.3
R13376 VSS.n5387 VSS.n5386 9.3
R13377 VSS.n5393 VSS.n5392 9.3
R13378 VSS.n5396 VSS.n5395 9.3
R13379 VSS.n5396 VSS.n5236 9.3
R13380 VSS.n5241 VSS.n5236 9.3
R13381 VSS.n5408 VSS.n5407 9.3
R13382 VSS.n5405 VSS.n5404 9.3
R13383 VSS.n5404 VSS.n5403 9.3
R13384 VSS.n5403 VSS.n5402 9.3
R13385 VSS.n5230 VSS.n1524 9.3
R13386 VSS.n5227 VSS.n1530 9.3
R13387 VSS.n1530 VSS.n1529 9.3
R13388 VSS.n1529 VSS.n1528 9.3
R13389 VSS.n5226 VSS.n5225 9.3
R13390 VSS.n5216 VSS.n5215 9.3
R13391 VSS.n5216 VSS.n1534 9.3
R13392 VSS.n5220 VSS.n1534 9.3
R13393 VSS.n5214 VSS.n5213 9.3
R13394 VSS.n5211 VSS.n1541 9.3
R13395 VSS.n5211 VSS.n5210 9.3
R13396 VSS.n5210 VSS.n5209 9.3
R13397 VSS.n5204 VSS.n5203 9.3
R13398 VSS.n5201 VSS.n5200 9.3
R13399 VSS.n5200 VSS.n1544 9.3
R13400 VSS.n1544 VSS.n1543 9.3
R13401 VSS.n1552 VSS.n1546 9.3
R13402 VSS.n5193 VSS.n5192 9.3
R13403 VSS.n5194 VSS.n5193 9.3
R13404 VSS.n5195 VSS.n5194 9.3
R13405 VSS.n5190 VSS.n5189 9.3
R13406 VSS.n5181 VSS.n5180 9.3
R13407 VSS.n5181 VSS.n1556 9.3
R13408 VSS.n5185 VSS.n1556 9.3
R13409 VSS.n5179 VSS.n5178 9.3
R13410 VSS.n5176 VSS.n1562 9.3
R13411 VSS.n5176 VSS.n5175 9.3
R13412 VSS.n5175 VSS.n5174 9.3
R13413 VSS.n5169 VSS.n5168 9.3
R13414 VSS.n5166 VSS.n5165 9.3
R13415 VSS.n5165 VSS.n1565 9.3
R13416 VSS.n1565 VSS.n1564 9.3
R13417 VSS.n1573 VSS.n1567 9.3
R13418 VSS.n5158 VSS.n5157 9.3
R13419 VSS.n5159 VSS.n5158 9.3
R13420 VSS.n5160 VSS.n5159 9.3
R13421 VSS.n5155 VSS.n5154 9.3
R13422 VSS.n5146 VSS.n5145 9.3
R13423 VSS.n5146 VSS.n1577 9.3
R13424 VSS.n5150 VSS.n1577 9.3
R13425 VSS.n5144 VSS.n5143 9.3
R13426 VSS.n5141 VSS.n1583 9.3
R13427 VSS.n5141 VSS.n5140 9.3
R13428 VSS.n5140 VSS.n5139 9.3
R13429 VSS.n1172 VSS.n1089 9.3
R13430 VSS.n1173 VSS.n1172 9.3
R13431 VSS.n1174 VSS.n1173 9.3
R13432 VSS.n1169 VSS.n1094 9.3
R13433 VSS.n6708 VSS.n6707 9.3
R13434 VSS.n6707 VSS.n6607 9.3
R13435 VSS.n6710 VSS.n6709 9.3
R13436 VSS.n6714 VSS.n6713 9.3
R13437 VSS.n6713 VSS.n6712 9.3
R13438 VSS.n6720 VSS.n6719 9.3
R13439 VSS.n6719 VSS.n6718 9.3
R13440 VSS.n6722 VSS.n6721 9.3
R13441 VSS.n6726 VSS.n6725 9.3
R13442 VSS.n6725 VSS.n6724 9.3
R13443 VSS.n6732 VSS.n6731 9.3
R13444 VSS.n6731 VSS.n6730 9.3
R13445 VSS.n6733 VSS.n6678 9.3
R13446 VSS.n6737 VSS.n6677 9.3
R13447 VSS.n6737 VSS.n6736 9.3
R13448 VSS.n6746 VSS.n6744 9.3
R13449 VSS.n6746 VSS.n6745 9.3
R13450 VSS.n6676 VSS.n6618 9.3
R13451 VSS.n6673 VSS.n6620 9.3
R13452 VSS.n6673 VSS.n6617 9.3
R13453 VSS.n6705 VSS.n6704 9.3
R13454 VSS.n6716 VSS.n6715 9.3
R13455 VSS.n6728 VSS.n6727 9.3
R13456 VSS.n6742 VSS.n6741 9.3
R13457 VSS.n6703 VSS.n6702 9.3
R13458 VSS.n6702 VSS.n6582 9.3
R13459 VSS.n6580 VSS.n6579 9.3
R13460 VSS.n6798 VSS.n6797 9.3
R13461 VSS.n6797 VSS.n6517 9.3
R13462 VSS.n6800 VSS.n6799 9.3
R13463 VSS.n6804 VSS.n6803 9.3
R13464 VSS.n6803 VSS.n6802 9.3
R13465 VSS.n6810 VSS.n6809 9.3
R13466 VSS.n6809 VSS.n6808 9.3
R13467 VSS.n6812 VSS.n6811 9.3
R13468 VSS.n6816 VSS.n6815 9.3
R13469 VSS.n6815 VSS.n6814 9.3
R13470 VSS.n6822 VSS.n6821 9.3
R13471 VSS.n6821 VSS.n6820 9.3
R13472 VSS.n6823 VSS.n6768 9.3
R13473 VSS.n6827 VSS.n6767 9.3
R13474 VSS.n6827 VSS.n6826 9.3
R13475 VSS.n6836 VSS.n6834 9.3
R13476 VSS.n6836 VSS.n6835 9.3
R13477 VSS.n6766 VSS.n6528 9.3
R13478 VSS.n6763 VSS.n6530 9.3
R13479 VSS.n6763 VSS.n6527 9.3
R13480 VSS.n6795 VSS.n6794 9.3
R13481 VSS.n6806 VSS.n6805 9.3
R13482 VSS.n6818 VSS.n6817 9.3
R13483 VSS.n6832 VSS.n6831 9.3
R13484 VSS.n6793 VSS.n6792 9.3
R13485 VSS.n6792 VSS.n6492 9.3
R13486 VSS.n6490 VSS.n6489 9.3
R13487 VSS.n6888 VSS.n6887 9.3
R13488 VSS.n6887 VSS.n6427 9.3
R13489 VSS.n6890 VSS.n6889 9.3
R13490 VSS.n6894 VSS.n6893 9.3
R13491 VSS.n6893 VSS.n6892 9.3
R13492 VSS.n6900 VSS.n6899 9.3
R13493 VSS.n6899 VSS.n6898 9.3
R13494 VSS.n6902 VSS.n6901 9.3
R13495 VSS.n6906 VSS.n6905 9.3
R13496 VSS.n6905 VSS.n6904 9.3
R13497 VSS.n6912 VSS.n6911 9.3
R13498 VSS.n6911 VSS.n6910 9.3
R13499 VSS.n6913 VSS.n6858 9.3
R13500 VSS.n6917 VSS.n6857 9.3
R13501 VSS.n6917 VSS.n6916 9.3
R13502 VSS.n6926 VSS.n6924 9.3
R13503 VSS.n6926 VSS.n6925 9.3
R13504 VSS.n6856 VSS.n6438 9.3
R13505 VSS.n6853 VSS.n6440 9.3
R13506 VSS.n6853 VSS.n6437 9.3
R13507 VSS.n6885 VSS.n6884 9.3
R13508 VSS.n6896 VSS.n6895 9.3
R13509 VSS.n6908 VSS.n6907 9.3
R13510 VSS.n6922 VSS.n6921 9.3
R13511 VSS.n6883 VSS.n6882 9.3
R13512 VSS.n6882 VSS.n6402 9.3
R13513 VSS.n6400 VSS.n6399 9.3
R13514 VSS.n5840 VSS.n5838 9.3
R13515 VSS.n6370 VSS.n6369 9.3
R13516 VSS.n6306 VSS.n6305 9.3
R13517 VSS.n6242 VSS.n6241 9.3
R13518 VSS.n6245 VSS.n6244 9.3
R13519 VSS.n6246 VSS.n6245 9.3
R13520 VSS.n6175 VSS.n6173 9.3
R13521 VSS.n6175 VSS.n6174 9.3
R13522 VSS.n6159 VSS.n6157 9.3
R13523 VSS.n6159 VSS.n6158 9.3
R13524 VSS.n6143 VSS.n6141 9.3
R13525 VSS.n6143 VSS.n6142 9.3
R13526 VSS.n6127 VSS.n6073 9.3
R13527 VSS.n6127 VSS.n6126 9.3
R13528 VSS.n6132 VSS.n6131 9.3
R13529 VSS.n6135 VSS.n6133 9.3
R13530 VSS.n6135 VSS.n6134 9.3
R13531 VSS.n6140 VSS.n6139 9.3
R13532 VSS.n6148 VSS.n6147 9.3
R13533 VSS.n6151 VSS.n6149 9.3
R13534 VSS.n6151 VSS.n6150 9.3
R13535 VSS.n6156 VSS.n6155 9.3
R13536 VSS.n6164 VSS.n6163 9.3
R13537 VSS.n6167 VSS.n6165 9.3
R13538 VSS.n6167 VSS.n6166 9.3
R13539 VSS.n6172 VSS.n6171 9.3
R13540 VSS.n6180 VSS.n6179 9.3
R13541 VSS.n6183 VSS.n6181 9.3
R13542 VSS.n6183 VSS.n6182 9.3
R13543 VSS.n6188 VSS.n6187 9.3
R13544 VSS.n6309 VSS.n6308 9.3
R13545 VSS.n6310 VSS.n6309 9.3
R13546 VSS.n6059 VSS.n6057 9.3
R13547 VSS.n6059 VSS.n6058 9.3
R13548 VSS.n6043 VSS.n6041 9.3
R13549 VSS.n6043 VSS.n6042 9.3
R13550 VSS.n6027 VSS.n6025 9.3
R13551 VSS.n6027 VSS.n6026 9.3
R13552 VSS.n6011 VSS.n5957 9.3
R13553 VSS.n6011 VSS.n6010 9.3
R13554 VSS.n6016 VSS.n6015 9.3
R13555 VSS.n6019 VSS.n6017 9.3
R13556 VSS.n6019 VSS.n6018 9.3
R13557 VSS.n6024 VSS.n6023 9.3
R13558 VSS.n6032 VSS.n6031 9.3
R13559 VSS.n6035 VSS.n6033 9.3
R13560 VSS.n6035 VSS.n6034 9.3
R13561 VSS.n6040 VSS.n6039 9.3
R13562 VSS.n6048 VSS.n6047 9.3
R13563 VSS.n6051 VSS.n6049 9.3
R13564 VSS.n6051 VSS.n6050 9.3
R13565 VSS.n6056 VSS.n6055 9.3
R13566 VSS.n6064 VSS.n6063 9.3
R13567 VSS.n6067 VSS.n6065 9.3
R13568 VSS.n6067 VSS.n6066 9.3
R13569 VSS.n6072 VSS.n6071 9.3
R13570 VSS.n6373 VSS.n6372 9.3
R13571 VSS.n6374 VSS.n6373 9.3
R13572 VSS.n5943 VSS.n5941 9.3
R13573 VSS.n5943 VSS.n5942 9.3
R13574 VSS.n5927 VSS.n5925 9.3
R13575 VSS.n5927 VSS.n5926 9.3
R13576 VSS.n5911 VSS.n5909 9.3
R13577 VSS.n5911 VSS.n5910 9.3
R13578 VSS.n5895 VSS.n5841 9.3
R13579 VSS.n5895 VSS.n5894 9.3
R13580 VSS.n5900 VSS.n5899 9.3
R13581 VSS.n5903 VSS.n5901 9.3
R13582 VSS.n5903 VSS.n5902 9.3
R13583 VSS.n5908 VSS.n5907 9.3
R13584 VSS.n5916 VSS.n5915 9.3
R13585 VSS.n5919 VSS.n5917 9.3
R13586 VSS.n5919 VSS.n5918 9.3
R13587 VSS.n5924 VSS.n5923 9.3
R13588 VSS.n5932 VSS.n5931 9.3
R13589 VSS.n5935 VSS.n5933 9.3
R13590 VSS.n5935 VSS.n5934 9.3
R13591 VSS.n5940 VSS.n5939 9.3
R13592 VSS.n5948 VSS.n5947 9.3
R13593 VSS.n5951 VSS.n5949 9.3
R13594 VSS.n5951 VSS.n5950 9.3
R13595 VSS.n5956 VSS.n5955 9.3
R13596 VSS.n6995 VSS.n5836 9.3
R13597 VSS.n6995 VSS.n6994 9.3
R13598 VSS.n7007 VSS.n5824 9.3
R13599 VSS.n7007 VSS.n7006 9.3
R13600 VSS.n7019 VSS.n5812 9.3
R13601 VSS.n7019 VSS.n7018 9.3
R13602 VSS.n7031 VSS.n5800 9.3
R13603 VSS.n7031 VSS.n7030 9.3
R13604 VSS.n7044 VSS.n7043 9.3
R13605 VSS.n7043 VSS.n7042 9.3
R13606 VSS.n5793 VSS.n5791 9.3
R13607 VSS.n7037 VSS.n5794 9.3
R13608 VSS.n7037 VSS.n7036 9.3
R13609 VSS.n5799 VSS.n5796 9.3
R13610 VSS.n5805 VSS.n5802 9.3
R13611 VSS.n7025 VSS.n5806 9.3
R13612 VSS.n7025 VSS.n7024 9.3
R13613 VSS.n5811 VSS.n5808 9.3
R13614 VSS.n5816 VSS.n5814 9.3
R13615 VSS.n7013 VSS.n5817 9.3
R13616 VSS.n7013 VSS.n7012 9.3
R13617 VSS.n5823 VSS.n5819 9.3
R13618 VSS.n5829 VSS.n5826 9.3
R13619 VSS.n7001 VSS.n5830 9.3
R13620 VSS.n7001 VSS.n7000 9.3
R13621 VSS.n5835 VSS.n5832 9.3
R13622 VSS.n381 VSS.n380 9.3
R13623 VSS.n380 VSS.n379 9.3
R13624 VSS.n370 VSS.n369 9.3
R13625 VSS.n365 VSS.n364 9.3
R13626 VSS.n401 VSS.n400 9.3
R13627 VSS.n356 VSS.n355 9.3
R13628 VSS.n352 VSS.n351 9.3
R13629 VSS.n347 VSS.n346 9.3
R13630 VSS.n383 VSS.n382 9.3
R13631 VSS.n388 VSS.n387 9.3
R13632 VSS.n387 VSS.n386 9.3
R13633 VSS.n390 VSS.n389 9.3
R13634 VSS.n398 VSS.n397 9.3
R13635 VSS.n397 VSS.n396 9.3
R13636 VSS.n399 VSS.n363 9.3
R13637 VSS.n402 VSS.n359 9.3
R13638 VSS.n402 VSS.n362 9.3
R13639 VSS.n411 VSS.n410 9.3
R13640 VSS.n412 VSS.n411 9.3
R13641 VSS.n416 VSS.n415 9.3
R13642 VSS.n418 VSS.n417 9.3
R13643 VSS.n419 VSS.n418 9.3
R13644 VSS.n423 VSS.n422 9.3
R13645 VSS.n425 VSS.n424 9.3
R13646 VSS.n426 VSS.n425 9.3
R13647 VSS.n431 VSS.n430 9.3
R13648 VSS.n432 VSS.n345 9.3
R13649 VSS.n345 VSS.n344 9.3
R13650 VSS.n435 VSS.n343 9.3
R13651 VSS.n434 VSS.n433 9.3
R13652 VSS.n374 VSS.n373 9.3
R13653 VSS.n377 VSS.n376 9.3
R13654 VSS.n18019 VSS.n18018 9.3
R13655 VSS.n18226 VSS.n18136 9.3
R13656 VSS.n18218 VSS.n18140 9.3
R13657 VSS.n18209 VSS.n18146 9.3
R13658 VSS.n18148 VSS.n18147 9.3
R13659 VSS.n18193 VSS.n18192 9.3
R13660 VSS.n18157 VSS.n18156 9.3
R13661 VSS.n18162 VSS.n18161 9.3
R13662 VSS.n18166 VSS.n18165 9.3
R13663 VSS.n18169 VSS.n18168 9.3
R13664 VSS.n18173 VSS.n18172 9.3
R13665 VSS.n18172 VSS.n18171 9.3
R13666 VSS.n18175 VSS.n18174 9.3
R13667 VSS.n18180 VSS.n18179 9.3
R13668 VSS.n18179 VSS.n18178 9.3
R13669 VSS.n18182 VSS.n18181 9.3
R13670 VSS.n18190 VSS.n18189 9.3
R13671 VSS.n18189 VSS.n18188 9.3
R13672 VSS.n18191 VSS.n18155 9.3
R13673 VSS.n18194 VSS.n18151 9.3
R13674 VSS.n18194 VSS.n18154 9.3
R13675 VSS.n18203 VSS.n18202 9.3
R13676 VSS.n18204 VSS.n18203 9.3
R13677 VSS.n18208 VSS.n18207 9.3
R13678 VSS.n18211 VSS.n18210 9.3
R13679 VSS.n18212 VSS.n18211 9.3
R13680 VSS.n18145 VSS.n18141 9.3
R13681 VSS.n18217 VSS.n18216 9.3
R13682 VSS.n18216 VSS.n18139 9.3
R13683 VSS.n18220 VSS.n18219 9.3
R13684 VSS.n18225 VSS.n18138 9.3
R13685 VSS.n18225 VSS.n18224 9.3
R13686 VSS.n18228 VSS.n18227 9.3
R13687 VSS.n2377 VSS.n2375 9.066
R13688 VSS.n2467 VSS.n2465 9.066
R13689 VSS.n2557 VSS.n2555 9.066
R13690 VSS.n2647 VSS.n2645 9.066
R13691 VSS.n2737 VSS.n2735 9.066
R13692 VSS.n2827 VSS.n2825 9.066
R13693 VSS.n2917 VSS.n2915 9.066
R13694 VSS.n3007 VSS.n3005 9.066
R13695 VSS.n6251 VSS.n6250 9.066
R13696 VSS.n6315 VSS.n6314 9.066
R13697 VSS.n6379 VSS.n6378 9.066
R13698 VSS.n6940 VSS.n6939 9.066
R13699 VSS.n6850 VSS.n6849 9.066
R13700 VSS.n6760 VSS.n6759 9.066
R13701 VSS.n6670 VSS.n6669 9.066
R13702 VSS.n1166 VSS.n1094 8.921
R13703 VSS.n4836 VSS.n3096 8.921
R13704 VSS.n408 VSS.n407 8.855
R13705 VSS.n18200 VSS.n18199 8.855
R13706 VSS VSS.n18089 8.809
R13707 VSS.n17881 VSS.n17880 8.791
R13708 VSS.n18232 VSS 8.735
R13709 VSS.n14642 VSS.n14641 8.533
R13710 VSS.n16570 VSS.n16569 8.533
R13711 VSS.n10691 VSS.n10690 8.533
R13712 VSS.n12619 VSS.n12618 8.533
R13713 VSS.n7259 VSS.n7258 8.533
R13714 VSS.n9187 VSS.n9186 8.533
R13715 VSS.n1654 VSS.n1652 8.533
R13716 VSS.n1167 VSS.n1165 8.533
R13717 VSS.n3814 VSS.n3446 8.533
R13718 VSS.n5129 VSS.n5128 8.533
R13719 VSS.n17809 VSS.n17805 8.533
R13720 VSS.n10578 VSS.n10566 8.454
R13721 VSS.n396 VSS.n395 8.275
R13722 VSS.n419 VSS.n353 8.275
R13723 VSS.n18188 VSS.n18187 8.275
R13724 VSS.n18212 VSS.n18143 8.275
R13725 VSS VSS.n17610 8.265
R13726 VSS.n14279 VSS.n14278 8.156
R13727 VSS.n14459 VSS.n14458 8.156
R13728 VSS.n12796 VSS.n12795 8.156
R13729 VSS.n12976 VSS.n12975 8.156
R13730 VSS.n13156 VSS.n13155 8.156
R13731 VSS.n13336 VSS.n13335 8.156
R13732 VSS.n13516 VSS.n13515 8.156
R13733 VSS.n13696 VSS.n13695 8.156
R13734 VSS.n13876 VSS.n13875 8.156
R13735 VSS.n14056 VSS.n14055 8.156
R13736 VSS.n6752 VSS.n6751 8.156
R13737 VSS.n6842 VSS.n6841 8.156
R13738 VSS.n6932 VSS.n6931 8.156
R13739 VSS.n438 VSS.n437 8.147
R13740 VSS.n5135 VSS.n5134 8.145
R13741 VSS.n3808 VSS.n3451 8.145
R13742 VSS.n7059 VSS.n7047 8.133
R13743 VSS.n17610 VSS.n17609 7.548
R13744 VSS.n17531 VSS.n17530 7.464
R13745 VSS.n17363 VSS.n17362 7.464
R13746 VSS.n17195 VSS.n17194 7.464
R13747 VSS.n17027 VSS.n17026 7.464
R13748 VSS.n16859 VSS.n16858 7.464
R13749 VSS.n16691 VSS.n16690 7.464
R13750 VSS.n10496 VSS.n10495 7.464
R13751 VSS.n6249 VSS.n6248 7.464
R13752 VSS.n6313 VSS.n6312 7.464
R13753 VSS.n6377 VSS.n6376 7.464
R13754 VSS.n6942 VSS.n6941 7.464
R13755 VSS.t64 VSS.n6247 7.262
R13756 VSS.t76 VSS.n6311 7.262
R13757 VSS.t74 VSS.n6375 7.262
R13758 VSS.n5837 VSS.t68 7.262
R13759 VSS.n16464 VSS.n16463 7.24
R13760 VSS.n16208 VSS.n16207 7.24
R13761 VSS.n15964 VSS.n15963 7.24
R13762 VSS.n15720 VSS.n15719 7.24
R13763 VSS.n15476 VSS.n15475 7.24
R13764 VSS.n15232 VSS.n15231 7.24
R13765 VSS.n14988 VSS.n14987 7.24
R13766 VSS.n14732 VSS.n14731 7.24
R13767 VSS.n12513 VSS.n12512 7.24
R13768 VSS.n12257 VSS.n12256 7.24
R13769 VSS.n12013 VSS.n12012 7.24
R13770 VSS.n11769 VSS.n11768 7.24
R13771 VSS.n11525 VSS.n11524 7.24
R13772 VSS.n11281 VSS.n11280 7.24
R13773 VSS.n11037 VSS.n11036 7.24
R13774 VSS.n10781 VSS.n10780 7.24
R13775 VSS.n9081 VSS.n9080 7.24
R13776 VSS.n8825 VSS.n8824 7.24
R13777 VSS.n8581 VSS.n8580 7.24
R13778 VSS.n8337 VSS.n8336 7.24
R13779 VSS.n8093 VSS.n8092 7.24
R13780 VSS.n7849 VSS.n7848 7.24
R13781 VSS.n7605 VSS.n7604 7.24
R13782 VSS.n7349 VSS.n7348 7.24
R13783 VSS.n1030 VSS.n1028 7.24
R13784 VSS.n1248 VSS.n1247 7.24
R13785 VSS.n1039 VSS.n1037 7.24
R13786 VSS.n1049 VSS.n1047 7.24
R13787 VSS.n1225 VSS.n1224 7.24
R13788 VSS.n1058 VSS.n1056 7.24
R13789 VSS.n1068 VSS.n1066 7.24
R13790 VSS.n1202 VSS.n1201 7.24
R13791 VSS.n1077 VSS.n1075 7.24
R13792 VSS.n1087 VSS.n1085 7.24
R13793 VSS.n1179 VSS.n1178 7.24
R13794 VSS.n927 VSS.n926 7.24
R13795 VSS.n935 VSS.n704 7.24
R13796 VSS.n946 VSS.n945 7.24
R13797 VSS.n697 VSS.n692 7.24
R13798 VSS.n962 VSS.n961 7.24
R13799 VSS.n970 VSS.n683 7.24
R13800 VSS.n981 VSS.n980 7.24
R13801 VSS.n676 VSS.n671 7.24
R13802 VSS.n997 VSS.n996 7.24
R13803 VSS.n1005 VSS.n662 7.24
R13804 VSS.n1016 VSS.n1015 7.24
R13805 VSS.n788 VSS.n776 7.24
R13806 VSS.n799 VSS.n798 7.24
R13807 VSS.n769 VSS.n764 7.24
R13808 VSS.n815 VSS.n814 7.24
R13809 VSS.n823 VSS.n755 7.24
R13810 VSS.n834 VSS.n833 7.24
R13811 VSS.n748 VSS.n743 7.24
R13812 VSS.n850 VSS.n849 7.24
R13813 VSS.n858 VSS.n734 7.24
R13814 VSS.n869 VSS.n868 7.24
R13815 VSS.n727 VSS.n726 7.24
R13816 VSS.n5600 VSS.n5599 7.24
R13817 VSS.n530 VSS.n528 7.24
R13818 VSS.n5771 VSS.n5770 7.24
R13819 VSS.n539 VSS.n537 7.24
R13820 VSS.n549 VSS.n547 7.24
R13821 VSS.n5748 VSS.n5747 7.24
R13822 VSS.n558 VSS.n556 7.24
R13823 VSS.n568 VSS.n566 7.24
R13824 VSS.n5725 VSS.n5724 7.24
R13825 VSS.n577 VSS.n575 7.24
R13826 VSS.n587 VSS.n585 7.24
R13827 VSS.n5502 VSS.n1439 7.24
R13828 VSS.n5513 VSS.n5512 7.24
R13829 VSS.n1432 VSS.n1427 7.24
R13830 VSS.n5529 VSS.n5528 7.24
R13831 VSS.n5537 VSS.n1418 7.24
R13832 VSS.n5548 VSS.n5547 7.24
R13833 VSS.n1411 VSS.n1406 7.24
R13834 VSS.n5564 VSS.n5563 7.24
R13835 VSS.n5572 VSS.n1397 7.24
R13836 VSS.n5584 VSS.n5583 7.24
R13837 VSS.n5590 VSS.n5589 7.24
R13838 VSS.n5392 VSS.n5391 7.24
R13839 VSS.n5246 VSS.n5244 7.24
R13840 VSS.n5256 VSS.n5254 7.24
R13841 VSS.n5369 VSS.n5368 7.24
R13842 VSS.n5265 VSS.n5263 7.24
R13843 VSS.n5275 VSS.n5273 7.24
R13844 VSS.n5346 VSS.n5345 7.24
R13845 VSS.n5284 VSS.n5282 7.24
R13846 VSS.n5294 VSS.n5292 7.24
R13847 VSS.n5323 VSS.n5322 7.24
R13848 VSS.n5304 VSS.n5301 7.24
R13849 VSS.n5143 VSS.n1580 7.24
R13850 VSS.n5154 VSS.n5153 7.24
R13851 VSS.n1573 VSS.n1568 7.24
R13852 VSS.n5170 VSS.n5169 7.24
R13853 VSS.n5178 VSS.n1559 7.24
R13854 VSS.n5189 VSS.n5188 7.24
R13855 VSS.n1552 VSS.n1547 7.24
R13856 VSS.n5205 VSS.n5204 7.24
R13857 VSS.n5213 VSS.n1538 7.24
R13858 VSS.n5225 VSS.n5224 7.24
R13859 VSS.n5231 VSS.n5230 7.24
R13860 VSS.n4774 VSS.n4772 7.24
R13861 VSS.n4915 VSS.n4914 7.24
R13862 VSS.n4783 VSS.n4781 7.24
R13863 VSS.n4793 VSS.n4791 7.24
R13864 VSS.n4892 VSS.n4891 7.24
R13865 VSS.n4802 VSS.n4800 7.24
R13866 VSS.n4812 VSS.n4810 7.24
R13867 VSS.n4869 VSS.n4868 7.24
R13868 VSS.n4821 VSS.n4819 7.24
R13869 VSS.n4831 VSS.n4829 7.24
R13870 VSS.n4846 VSS.n4845 7.24
R13871 VSS.n4662 VSS.n4660 7.24
R13872 VSS.n5008 VSS.n5007 7.24
R13873 VSS.n4671 VSS.n4669 7.24
R13874 VSS.n4681 VSS.n4679 7.24
R13875 VSS.n4985 VSS.n4984 7.24
R13876 VSS.n4690 VSS.n4688 7.24
R13877 VSS.n4700 VSS.n4698 7.24
R13878 VSS.n4962 VSS.n4961 7.24
R13879 VSS.n4709 VSS.n4707 7.24
R13880 VSS.n4719 VSS.n4717 7.24
R13881 VSS.n4939 VSS.n4938 7.24
R13882 VSS.n4554 VSS.n4553 7.24
R13883 VSS.n3211 VSS.n3206 7.24
R13884 VSS.n4570 VSS.n4569 7.24
R13885 VSS.n4578 VSS.n3197 7.24
R13886 VSS.n4589 VSS.n4588 7.24
R13887 VSS.n3190 VSS.n3185 7.24
R13888 VSS.n4605 VSS.n4604 7.24
R13889 VSS.n4613 VSS.n3176 7.24
R13890 VSS.n4624 VSS.n4623 7.24
R13891 VSS.n3169 VSS.n3164 7.24
R13892 VSS.n4640 VSS.n4639 7.24
R13893 VSS.n4184 VSS.n4182 7.24
R13894 VSS.n4306 VSS.n4305 7.24
R13895 VSS.n4193 VSS.n4191 7.24
R13896 VSS.n4203 VSS.n4201 7.24
R13897 VSS.n4283 VSS.n4282 7.24
R13898 VSS.n4212 VSS.n4210 7.24
R13899 VSS.n4222 VSS.n4220 7.24
R13900 VSS.n4260 VSS.n4259 7.24
R13901 VSS.n4231 VSS.n4229 7.24
R13902 VSS.n4238 VSS.n4237 7.24
R13903 VSS.n4537 VSS.n4536 7.24
R13904 VSS.n4072 VSS.n4070 7.24
R13905 VSS.n4399 VSS.n4398 7.24
R13906 VSS.n4081 VSS.n4079 7.24
R13907 VSS.n4091 VSS.n4089 7.24
R13908 VSS.n4376 VSS.n4375 7.24
R13909 VSS.n4100 VSS.n4098 7.24
R13910 VSS.n4110 VSS.n4108 7.24
R13911 VSS.n4353 VSS.n4352 7.24
R13912 VSS.n4119 VSS.n4117 7.24
R13913 VSS.n4129 VSS.n4127 7.24
R13914 VSS.n4330 VSS.n4329 7.24
R13915 VSS.n3969 VSS.n3968 7.24
R13916 VSS.n3977 VSS.n3374 7.24
R13917 VSS.n3988 VSS.n3987 7.24
R13918 VSS.n3367 VSS.n3362 7.24
R13919 VSS.n4004 VSS.n4003 7.24
R13920 VSS.n4012 VSS.n3353 7.24
R13921 VSS.n4023 VSS.n4022 7.24
R13922 VSS.n3346 VSS.n3341 7.24
R13923 VSS.n4039 VSS.n4038 7.24
R13924 VSS.n4047 VSS.n3332 7.24
R13925 VSS.n4058 VSS.n4057 7.24
R13926 VSS.n3572 VSS.n3570 7.24
R13927 VSS.n3702 VSS.n3701 7.24
R13928 VSS.n3581 VSS.n3579 7.24
R13929 VSS.n3591 VSS.n3589 7.24
R13930 VSS.n3679 VSS.n3678 7.24
R13931 VSS.n3600 VSS.n3598 7.24
R13932 VSS.n3610 VSS.n3608 7.24
R13933 VSS.n3656 VSS.n3655 7.24
R13934 VSS.n3619 VSS.n3617 7.24
R13935 VSS.n3633 VSS.n3627 7.24
R13936 VSS.n3631 VSS.n3630 7.24
R13937 VSS.n3460 VSS.n3457 7.24
R13938 VSS.n3795 VSS.n3794 7.24
R13939 VSS.n3469 VSS.n3467 7.24
R13940 VSS.n3479 VSS.n3477 7.24
R13941 VSS.n3772 VSS.n3771 7.24
R13942 VSS.n3488 VSS.n3486 7.24
R13943 VSS.n3498 VSS.n3496 7.24
R13944 VSS.n3749 VSS.n3748 7.24
R13945 VSS.n3507 VSS.n3505 7.24
R13946 VSS.n3517 VSS.n3515 7.24
R13947 VSS.n3726 VSS.n3725 7.24
R13948 VSS.n14311 VSS.n14310 7.111
R13949 VSS.n14132 VSS.n14131 7.111
R13950 VSS.n17596 VSS.n17595 7.111
R13951 VSS.n17428 VSS.n17427 7.111
R13952 VSS.n17260 VSS.n17259 7.111
R13953 VSS.n17092 VSS.n17091 7.111
R13954 VSS.n16924 VSS.n16923 7.111
R13955 VSS.n16756 VSS.n16755 7.111
R13956 VSS.n13908 VSS.n13907 7.111
R13957 VSS.n13728 VSS.n13727 7.111
R13958 VSS.n13548 VSS.n13547 7.111
R13959 VSS.n13368 VSS.n13367 7.111
R13960 VSS.n13188 VSS.n13187 7.111
R13961 VSS.n13008 VSS.n13007 7.111
R13962 VSS.n12828 VSS.n12827 7.111
R13963 VSS.n12649 VSS.n12648 7.111
R13964 VSS.n7168 VSS.n7167 7.111
R13965 VSS.n7156 VSS.n7155 7.111
R13966 VSS.n7144 VSS.n7143 7.111
R13967 VSS.n7132 VSS.n7131 7.111
R13968 VSS.n7120 VSS.n7119 7.111
R13969 VSS.n7108 VSS.n7107 7.111
R13970 VSS.n7096 VSS.n7095 7.111
R13971 VSS.n10563 VSS.n10561 7.111
R13972 VSS.n2375 VSS.n2374 7.111
R13973 VSS.n2465 VSS.n2284 7.111
R13974 VSS.n2555 VSS.n2194 7.111
R13975 VSS.n2645 VSS.n2104 7.111
R13976 VSS.n2735 VSS.n2014 7.111
R13977 VSS.n2825 VSS.n1924 7.111
R13978 VSS.n2915 VSS.n1834 7.111
R13979 VSS.n3005 VSS.n1744 7.111
R13980 VSS.n6251 VSS.n6074 7.111
R13981 VSS.n6315 VSS.n5958 7.111
R13982 VSS.n6379 VSS.n5842 7.111
R13983 VSS.n6945 VSS.n6939 7.111
R13984 VSS.n6849 VSS.n6488 7.111
R13985 VSS.n6759 VSS.n6578 7.111
R13986 VSS.n6669 VSS.n6668 7.111
R13987 VSS VSS.n17642 6.972
R13988 VSS VSS.n470 6.972
R13989 VSS.n18027 VSS 6.972
R13990 VSS.n14133 VSS.n14132 6.925
R13991 VSS.n12650 VSS.n12649 6.925
R13992 VSS.n2375 VSS.n2326 6.925
R13993 VSS.n6669 VSS.n6620 6.925
R13994 VSS.n14312 VSS.n14311 6.783
R13995 VSS.n17597 VSS.n17596 6.783
R13996 VSS.n17429 VSS.n17428 6.783
R13997 VSS.n17261 VSS.n17260 6.783
R13998 VSS.n17093 VSS.n17092 6.783
R13999 VSS.n16925 VSS.n16924 6.783
R14000 VSS.n16757 VSS.n16756 6.783
R14001 VSS.n13909 VSS.n13908 6.783
R14002 VSS.n13729 VSS.n13728 6.783
R14003 VSS.n13549 VSS.n13548 6.783
R14004 VSS.n13369 VSS.n13368 6.783
R14005 VSS.n13189 VSS.n13188 6.783
R14006 VSS.n13009 VSS.n13008 6.783
R14007 VSS.n12829 VSS.n12828 6.783
R14008 VSS.n9374 VSS.n7168 6.783
R14009 VSS.n9542 VSS.n7156 6.783
R14010 VSS.n9710 VSS.n7144 6.783
R14011 VSS.n9878 VSS.n7132 6.783
R14012 VSS.n10046 VSS.n7120 6.783
R14013 VSS.n10214 VSS.n7108 6.783
R14014 VSS.n10382 VSS.n7096 6.783
R14015 VSS.n2465 VSS.n2464 6.783
R14016 VSS.n2555 VSS.n2554 6.783
R14017 VSS.n2645 VSS.n2644 6.783
R14018 VSS.n2735 VSS.n2734 6.783
R14019 VSS.n2825 VSS.n2824 6.783
R14020 VSS.n2915 VSS.n2914 6.783
R14021 VSS.n3005 VSS.n3004 6.783
R14022 VSS.n6252 VSS.n6251 6.783
R14023 VSS.n6316 VSS.n6315 6.783
R14024 VSS.n6380 VSS.n6379 6.783
R14025 VSS.n6849 VSS.n6848 6.783
R14026 VSS.n6759 VSS.n6758 6.783
R14027 VSS.n16334 VSS.n16317 6.723
R14028 VSS.n16079 VSS.n16062 6.723
R14029 VSS.n15834 VSS.n15817 6.723
R14030 VSS.n15591 VSS.n15574 6.723
R14031 VSS.n15346 VSS.n15329 6.723
R14032 VSS.n15103 VSS.n15086 6.723
R14033 VSS.n14858 VSS.n14829 6.723
R14034 VSS.n12383 VSS.n12366 6.723
R14035 VSS.n12128 VSS.n12111 6.723
R14036 VSS.n11883 VSS.n11866 6.723
R14037 VSS.n11640 VSS.n11623 6.723
R14038 VSS.n11395 VSS.n11378 6.723
R14039 VSS.n11152 VSS.n11135 6.723
R14040 VSS.n10907 VSS.n10878 6.723
R14041 VSS.n8951 VSS.n8934 6.723
R14042 VSS.n8696 VSS.n8679 6.723
R14043 VSS.n8451 VSS.n8434 6.723
R14044 VSS.n8208 VSS.n8191 6.723
R14045 VSS.n7963 VSS.n7946 6.723
R14046 VSS.n7720 VSS.n7703 6.723
R14047 VSS.n7475 VSS.n7446 6.723
R14048 VSS.n1297 VSS.n637 6.723
R14049 VSS.n1322 VSS.n1321 6.723
R14050 VSS.n1348 VSS.n605 6.723
R14051 VSS.n5644 VSS.n1361 6.723
R14052 VSS.n1489 VSS.n1460 6.723
R14053 VSS.n5436 VSS.n1502 6.723
R14054 VSS.n5081 VSS.n5080 6.723
R14055 VSS.n5053 VSS.n3138 6.723
R14056 VSS.n3275 VSS.n3241 6.723
R14057 VSS.n4474 VSS.n3288 6.723
R14058 VSS.n4449 VSS.n4448 6.723
R14059 VSS.n3925 VSS.n3405 6.723
R14060 VSS.n3866 VSS.n3865 6.723
R14061 VSS VSS.n17769 6.216
R14062 VSS.n16334 VSS.n16333 6.206
R14063 VSS.n16079 VSS.n16078 6.206
R14064 VSS.n15834 VSS.n15833 6.206
R14065 VSS.n15591 VSS.n15590 6.206
R14066 VSS.n15346 VSS.n15345 6.206
R14067 VSS.n15103 VSS.n15102 6.206
R14068 VSS.n14858 VSS.n14857 6.206
R14069 VSS.n12383 VSS.n12382 6.206
R14070 VSS.n12128 VSS.n12127 6.206
R14071 VSS.n11883 VSS.n11882 6.206
R14072 VSS.n11640 VSS.n11639 6.206
R14073 VSS.n11395 VSS.n11394 6.206
R14074 VSS.n11152 VSS.n11151 6.206
R14075 VSS.n10907 VSS.n10906 6.206
R14076 VSS.n8951 VSS.n8950 6.206
R14077 VSS.n8696 VSS.n8695 6.206
R14078 VSS.n8451 VSS.n8450 6.206
R14079 VSS.n8208 VSS.n8207 6.206
R14080 VSS.n7963 VSS.n7962 6.206
R14081 VSS.n7720 VSS.n7719 6.206
R14082 VSS.n7475 VSS.n7474 6.206
R14083 VSS.n1298 VSS.n1297 6.206
R14084 VSS.n1322 VSS.n617 6.206
R14085 VSS.n5670 VSS.n605 6.206
R14086 VSS.n5645 VSS.n5644 6.206
R14087 VSS.n5462 VSS.n1460 6.206
R14088 VSS.n5437 VSS.n5436 6.206
R14089 VSS.n5080 VSS.n3123 6.206
R14090 VSS.n3253 VSS.n3138 6.206
R14091 VSS.n4500 VSS.n3241 6.206
R14092 VSS.n4474 VSS.n4473 6.206
R14093 VSS.n4448 VSS.n3307 6.206
R14094 VSS.n3925 VSS.n3924 6.206
R14095 VSS.n3865 VSS.n3419 6.206
R14096 VSS.n16571 VSS.n16570 6.201
R14097 VSS.n12620 VSS.n12619 6.201
R14098 VSS.n9188 VSS.n9187 6.201
R14099 VSS.n1168 VSS.n1167 6.201
R14100 VSS.n5130 VSS.n5129 6.201
R14101 VSS.n437 VSS.n436 6.156
R14102 VSS.n18229 VSS.n18135 6.084
R14103 VSS.n17921 VSS.n17920 6.076
R14104 VSS.n14083 VSS.n14082 5.903
R14105 VSS.n1021 VSS.n650 5.818
R14106 VSS.n885 VSS.n713 5.818
R14107 VSS.n5701 VSS.n590 5.818
R14108 VSS.n5617 VSS.n1380 5.818
R14109 VSS.n5494 VSS.n5493 5.818
R14110 VSS.n5409 VSS.n1521 5.818
R14111 VSS.n4766 VSS.n4760 5.818
R14112 VSS.n5022 VSS.n3155 5.818
R14113 VSS.n4543 VSS.n3218 5.818
R14114 VSS.n4176 VSS.n4170 5.818
R14115 VSS.n4063 VSS.n3320 5.818
R14116 VSS.n3951 VSS.n3383 5.818
R14117 VSS.n3564 VSS.n3558 5.818
R14118 VSS.n2315 VSS.n2309 5.655
R14119 VSS.n2376 VSS.n2315 5.655
R14120 VSS.n2225 VSS.n2219 5.655
R14121 VSS.n2466 VSS.n2225 5.655
R14122 VSS.n2135 VSS.n2129 5.655
R14123 VSS.n2556 VSS.n2135 5.655
R14124 VSS.n2045 VSS.n2039 5.655
R14125 VSS.n2646 VSS.n2045 5.655
R14126 VSS.n1955 VSS.n1949 5.655
R14127 VSS.n2736 VSS.n1955 5.655
R14128 VSS.n1865 VSS.n1859 5.655
R14129 VSS.n2826 VSS.n1865 5.655
R14130 VSS.n1775 VSS.n1769 5.655
R14131 VSS.n2916 VSS.n1775 5.655
R14132 VSS.n1685 VSS.n1679 5.655
R14133 VSS.n3006 VSS.n1685 5.655
R14134 VSS.n401 VSS.n363 5.647
R14135 VSS.n403 VSS.n360 5.647
R14136 VSS.n361 VSS.n358 5.647
R14137 VSS.n415 VSS.n356 5.647
R14138 VSS.n18193 VSS.n18155 5.647
R14139 VSS.n18195 VSS.n18152 5.647
R14140 VSS.n18153 VSS.n18150 5.647
R14141 VSS.n18207 VSS.n18148 5.647
R14142 VSS.n17921 VSS.n17770 5.559
R14143 VSS.n18018 VSS.n17924 5.464
R14144 VSS.n439 VSS.n331 5.454
R14145 VSS.n17579 VSS.t6 5.446
R14146 VSS.n17411 VSS.t2 5.446
R14147 VSS.n17243 VSS.t4 5.446
R14148 VSS.n17075 VSS.t12 5.446
R14149 VSS.n16907 VSS.t14 5.446
R14150 VSS.n16739 VSS.t0 5.446
R14151 VSS.n9367 VSS.n9366 5.446
R14152 VSS.n9535 VSS.n9534 5.446
R14153 VSS.n9703 VSS.n9702 5.446
R14154 VSS.n9871 VSS.n9870 5.446
R14155 VSS.n10039 VSS.n10038 5.446
R14156 VSS.n10207 VSS.n10206 5.446
R14157 VSS.n10375 VSS.n10374 5.446
R14158 VSS.n10543 VSS.t56 5.446
R14159 VSS.n2458 VSS.n2319 5.446
R14160 VSS.n2458 VSS.n2320 5.446
R14161 VSS.n2458 VSS.n2318 5.446
R14162 VSS.n2458 VSS.n2321 5.446
R14163 VSS.n2458 VSS.n2317 5.446
R14164 VSS.n2458 VSS.n2322 5.446
R14165 VSS.n2458 VSS.n2316 5.446
R14166 VSS.n2458 VSS.n2457 5.446
R14167 VSS.n2548 VSS.n2229 5.446
R14168 VSS.n2548 VSS.n2230 5.446
R14169 VSS.n2548 VSS.n2228 5.446
R14170 VSS.n2548 VSS.n2231 5.446
R14171 VSS.n2548 VSS.n2227 5.446
R14172 VSS.n2548 VSS.n2232 5.446
R14173 VSS.n2548 VSS.n2226 5.446
R14174 VSS.n2548 VSS.n2547 5.446
R14175 VSS.n2638 VSS.n2139 5.446
R14176 VSS.n2638 VSS.n2140 5.446
R14177 VSS.n2638 VSS.n2138 5.446
R14178 VSS.n2638 VSS.n2141 5.446
R14179 VSS.n2638 VSS.n2137 5.446
R14180 VSS.n2638 VSS.n2142 5.446
R14181 VSS.n2638 VSS.n2136 5.446
R14182 VSS.n2638 VSS.n2637 5.446
R14183 VSS.n2728 VSS.n2049 5.446
R14184 VSS.n2728 VSS.n2050 5.446
R14185 VSS.n2728 VSS.n2048 5.446
R14186 VSS.n2728 VSS.n2051 5.446
R14187 VSS.n2728 VSS.n2047 5.446
R14188 VSS.n2728 VSS.n2052 5.446
R14189 VSS.n2728 VSS.n2046 5.446
R14190 VSS.n2728 VSS.n2727 5.446
R14191 VSS.n2818 VSS.n1959 5.446
R14192 VSS.n2818 VSS.n1960 5.446
R14193 VSS.n2818 VSS.n1958 5.446
R14194 VSS.n2818 VSS.n1961 5.446
R14195 VSS.n2818 VSS.n1957 5.446
R14196 VSS.n2818 VSS.n1962 5.446
R14197 VSS.n2818 VSS.n1956 5.446
R14198 VSS.n2818 VSS.n2817 5.446
R14199 VSS.n2908 VSS.n1869 5.446
R14200 VSS.n2908 VSS.n1870 5.446
R14201 VSS.n2908 VSS.n1868 5.446
R14202 VSS.n2908 VSS.n1871 5.446
R14203 VSS.n2908 VSS.n1867 5.446
R14204 VSS.n2908 VSS.n1872 5.446
R14205 VSS.n2908 VSS.n1866 5.446
R14206 VSS.n2908 VSS.n2907 5.446
R14207 VSS.n2998 VSS.n1779 5.446
R14208 VSS.n2998 VSS.n1780 5.446
R14209 VSS.n2998 VSS.n1778 5.446
R14210 VSS.n2998 VSS.n1781 5.446
R14211 VSS.n2998 VSS.n1777 5.446
R14212 VSS.n2998 VSS.n1782 5.446
R14213 VSS.n2998 VSS.n1776 5.446
R14214 VSS.n2998 VSS.n2997 5.446
R14215 VSS.n3088 VSS.n1689 5.446
R14216 VSS.n3088 VSS.n1690 5.446
R14217 VSS.n3088 VSS.n1688 5.446
R14218 VSS.n3088 VSS.n1691 5.446
R14219 VSS.n3088 VSS.n1687 5.446
R14220 VSS.n3088 VSS.n1692 5.446
R14221 VSS.n3088 VSS.n1686 5.446
R14222 VSS.n3088 VSS.n3087 5.446
R14223 VSS.t64 VSS.n6102 5.446
R14224 VSS.t64 VSS.n6103 5.446
R14225 VSS.t64 VSS.n6101 5.446
R14226 VSS.t64 VSS.n6104 5.446
R14227 VSS.t64 VSS.n6105 5.446
R14228 VSS.t64 VSS.n6100 5.446
R14229 VSS.t64 VSS.n6106 5.446
R14230 VSS.t64 VSS.n6099 5.446
R14231 VSS.t76 VSS.n5986 5.446
R14232 VSS.t76 VSS.n5987 5.446
R14233 VSS.t76 VSS.n5985 5.446
R14234 VSS.t76 VSS.n5988 5.446
R14235 VSS.t76 VSS.n5989 5.446
R14236 VSS.t76 VSS.n5984 5.446
R14237 VSS.t76 VSS.n5990 5.446
R14238 VSS.t76 VSS.n5983 5.446
R14239 VSS.t74 VSS.n5870 5.446
R14240 VSS.t74 VSS.n5871 5.446
R14241 VSS.t74 VSS.n5869 5.446
R14242 VSS.t74 VSS.n5872 5.446
R14243 VSS.t74 VSS.n5873 5.446
R14244 VSS.t74 VSS.n5868 5.446
R14245 VSS.t74 VSS.n5874 5.446
R14246 VSS.t74 VSS.n5867 5.446
R14247 VSS.n6999 VSS.t68 5.446
R14248 VSS.n7011 VSS.t68 5.446
R14249 VSS.n7023 VSS.t68 5.446
R14250 VSS.n7035 VSS.t68 5.446
R14251 VSS.n7041 VSS.t68 5.446
R14252 VSS.n7029 VSS.t68 5.446
R14253 VSS.n7017 VSS.t68 5.446
R14254 VSS.n7005 VSS.t68 5.446
R14255 VSS.n6932 VSS.n6433 5.446
R14256 VSS.n6932 VSS.n6434 5.446
R14257 VSS.n6932 VSS.n6432 5.446
R14258 VSS.n6932 VSS.n6435 5.446
R14259 VSS.n6932 VSS.n6431 5.446
R14260 VSS.n6932 VSS.n6436 5.446
R14261 VSS.n6932 VSS.n6430 5.446
R14262 VSS.n6932 VSS.n6930 5.446
R14263 VSS.n6842 VSS.n6523 5.446
R14264 VSS.n6842 VSS.n6524 5.446
R14265 VSS.n6842 VSS.n6522 5.446
R14266 VSS.n6842 VSS.n6525 5.446
R14267 VSS.n6842 VSS.n6521 5.446
R14268 VSS.n6842 VSS.n6526 5.446
R14269 VSS.n6842 VSS.n6520 5.446
R14270 VSS.n6842 VSS.n6840 5.446
R14271 VSS.n6752 VSS.n6613 5.446
R14272 VSS.n6752 VSS.n6614 5.446
R14273 VSS.n6752 VSS.n6612 5.446
R14274 VSS.n6752 VSS.n6615 5.446
R14275 VSS.n6752 VSS.n6611 5.446
R14276 VSS.n6752 VSS.n6616 5.446
R14277 VSS.n6752 VSS.n6610 5.446
R14278 VSS.n6752 VSS.n6750 5.446
R14279 VSS.n7061 VSS 5.404
R14280 VSS.n498 VSS 5.404
R14281 VSS VSS.n17741 5.404
R14282 VSS VSS.n439 5.356
R14283 VSS VSS.n7059 5.337
R14284 VSS.n18018 VSS.n18017 5
R14285 VSS.n440 VSS 4.995
R14286 VSS.n390 VSS.n365 4.894
R14287 VSS.n393 VSS.n366 4.894
R14288 VSS.n414 VSS.n354 4.894
R14289 VSS.n422 VSS.n352 4.894
R14290 VSS.n18182 VSS.n18157 4.894
R14291 VSS.n18185 VSS.n18158 4.894
R14292 VSS.n18206 VSS.n18144 4.894
R14293 VSS.n18146 VSS.n18145 4.894
R14294 VSS.n10578 VSS.n10577 4.868
R14295 VSS.n14644 VSS.n14643 4.792
R14296 VSS.n10693 VSS.n10692 4.792
R14297 VSS.n7261 VSS.n7260 4.792
R14298 VSS.n3453 VSS.n3451 4.792
R14299 VSS.n7059 VSS 4.651
R14300 VSS.n16586 VSS.n16585 4.65
R14301 VSS.n14659 VSS.n14658 4.65
R14302 VSS.n14673 VSS.n14672 4.65
R14303 VSS.n14687 VSS.n14686 4.65
R14304 VSS.n14701 VSS.n14700 4.65
R14305 VSS.n14715 VSS.n14714 4.65
R14306 VSS.n14734 VSS.n14733 4.65
R14307 VSS.n14737 VSS.n14599 4.65
R14308 VSS.n14751 VSS.n14750 4.65
R14309 VSS.n14765 VSS.n14764 4.65
R14310 VSS.n14779 VSS.n14778 4.65
R14311 VSS.n14793 VSS.n14792 4.65
R14312 VSS.n14810 VSS.n14809 4.65
R14313 VSS.n14915 VSS.n14914 4.65
R14314 VSS.n14929 VSS.n14928 4.65
R14315 VSS.n14943 VSS.n14942 4.65
R14316 VSS.n14957 VSS.n14956 4.65
R14317 VSS.n14971 VSS.n14970 4.65
R14318 VSS.n14990 VSS.n14989 4.65
R14319 VSS.n14993 VSS.n14593 4.65
R14320 VSS.n15007 VSS.n15006 4.65
R14321 VSS.n15021 VSS.n15020 4.65
R14322 VSS.n15035 VSS.n15034 4.65
R14323 VSS.n15049 VSS.n15048 4.65
R14324 VSS.n15066 VSS.n15065 4.65
R14325 VSS.n15159 VSS.n15158 4.65
R14326 VSS.n15173 VSS.n15172 4.65
R14327 VSS.n15187 VSS.n15186 4.65
R14328 VSS.n15201 VSS.n15200 4.65
R14329 VSS.n15215 VSS.n15214 4.65
R14330 VSS.n15234 VSS.n15233 4.65
R14331 VSS.n15237 VSS.n14587 4.65
R14332 VSS.n15251 VSS.n15250 4.65
R14333 VSS.n15265 VSS.n15264 4.65
R14334 VSS.n15279 VSS.n15278 4.65
R14335 VSS.n15293 VSS.n15292 4.65
R14336 VSS.n15310 VSS.n15309 4.65
R14337 VSS.n15403 VSS.n15402 4.65
R14338 VSS.n15417 VSS.n15416 4.65
R14339 VSS.n15431 VSS.n15430 4.65
R14340 VSS.n15445 VSS.n15444 4.65
R14341 VSS.n15459 VSS.n15458 4.65
R14342 VSS.n15478 VSS.n15477 4.65
R14343 VSS.n15481 VSS.n14581 4.65
R14344 VSS.n15495 VSS.n15494 4.65
R14345 VSS.n15509 VSS.n15508 4.65
R14346 VSS.n15523 VSS.n15522 4.65
R14347 VSS.n15537 VSS.n15536 4.65
R14348 VSS.n15554 VSS.n15553 4.65
R14349 VSS.n15647 VSS.n15646 4.65
R14350 VSS.n15661 VSS.n15660 4.65
R14351 VSS.n15675 VSS.n15674 4.65
R14352 VSS.n15689 VSS.n15688 4.65
R14353 VSS.n15703 VSS.n15702 4.65
R14354 VSS.n15722 VSS.n15721 4.65
R14355 VSS.n15725 VSS.n14575 4.65
R14356 VSS.n15739 VSS.n15738 4.65
R14357 VSS.n15753 VSS.n15752 4.65
R14358 VSS.n15767 VSS.n15766 4.65
R14359 VSS.n15781 VSS.n15780 4.65
R14360 VSS.n15798 VSS.n15797 4.65
R14361 VSS.n15891 VSS.n15890 4.65
R14362 VSS.n15905 VSS.n15904 4.65
R14363 VSS.n15919 VSS.n15918 4.65
R14364 VSS.n15933 VSS.n15932 4.65
R14365 VSS.n15947 VSS.n15946 4.65
R14366 VSS.n15966 VSS.n15965 4.65
R14367 VSS.n15969 VSS.n14569 4.65
R14368 VSS.n15983 VSS.n15982 4.65
R14369 VSS.n15997 VSS.n15996 4.65
R14370 VSS.n16011 VSS.n16010 4.65
R14371 VSS.n16025 VSS.n16024 4.65
R14372 VSS.n16042 VSS.n16041 4.65
R14373 VSS.n16135 VSS.n16134 4.65
R14374 VSS.n16149 VSS.n16148 4.65
R14375 VSS.n16163 VSS.n16162 4.65
R14376 VSS.n16177 VSS.n16176 4.65
R14377 VSS.n16191 VSS.n16190 4.65
R14378 VSS.n16210 VSS.n16209 4.65
R14379 VSS.n16213 VSS.n14563 4.65
R14380 VSS.n16227 VSS.n16226 4.65
R14381 VSS.n16241 VSS.n16240 4.65
R14382 VSS.n16255 VSS.n16254 4.65
R14383 VSS.n16269 VSS.n16268 4.65
R14384 VSS.n16286 VSS.n16285 4.65
R14385 VSS.n16525 VSS.n16524 4.65
R14386 VSS.n16511 VSS.n16510 4.65
R14387 VSS.n16497 VSS.n16496 4.65
R14388 VSS.n16483 VSS.n16482 4.65
R14389 VSS.n16469 VSS.n14557 4.65
R14390 VSS.n16466 VSS.n16465 4.65
R14391 VSS.n16447 VSS.n16446 4.65
R14392 VSS.n16433 VSS.n16432 4.65
R14393 VSS.n16419 VSS.n16418 4.65
R14394 VSS.n16405 VSS.n16404 4.65
R14395 VSS.n16391 VSS.n16390 4.65
R14396 VSS.n16590 VSS.n14551 4.65
R14397 VSS.n16744 VSS.n16743 4.65
R14398 VSS.n16685 VSS.n16684 4.65
R14399 VSS.n16673 VSS.n16672 4.65
R14400 VSS.n16661 VSS.n16660 4.65
R14401 VSS.n16649 VSS.n16648 4.65
R14402 VSS.n16632 VSS.n16628 4.65
R14403 VSS.n16625 VSS.n16624 4.65
R14404 VSS.n16613 VSS.n16612 4.65
R14405 VSS.n16601 VSS.n16600 4.65
R14406 VSS.n16758 VSS.n14539 4.65
R14407 VSS.n16912 VSS.n16911 4.65
R14408 VSS.n16853 VSS.n16852 4.65
R14409 VSS.n16841 VSS.n16840 4.65
R14410 VSS.n16829 VSS.n16828 4.65
R14411 VSS.n16817 VSS.n16816 4.65
R14412 VSS.n16800 VSS.n16796 4.65
R14413 VSS.n16793 VSS.n16792 4.65
R14414 VSS.n16781 VSS.n16780 4.65
R14415 VSS.n16769 VSS.n16768 4.65
R14416 VSS.n16926 VSS.n14527 4.65
R14417 VSS.n17080 VSS.n17079 4.65
R14418 VSS.n17021 VSS.n17020 4.65
R14419 VSS.n17009 VSS.n17008 4.65
R14420 VSS.n16997 VSS.n16996 4.65
R14421 VSS.n16985 VSS.n16984 4.65
R14422 VSS.n16968 VSS.n16964 4.65
R14423 VSS.n16961 VSS.n16960 4.65
R14424 VSS.n16949 VSS.n16948 4.65
R14425 VSS.n16937 VSS.n16936 4.65
R14426 VSS.n17094 VSS.n14515 4.65
R14427 VSS.n17248 VSS.n17247 4.65
R14428 VSS.n17189 VSS.n17188 4.65
R14429 VSS.n17177 VSS.n17176 4.65
R14430 VSS.n17165 VSS.n17164 4.65
R14431 VSS.n17153 VSS.n17152 4.65
R14432 VSS.n17136 VSS.n17132 4.65
R14433 VSS.n17129 VSS.n17128 4.65
R14434 VSS.n17117 VSS.n17116 4.65
R14435 VSS.n17105 VSS.n17104 4.65
R14436 VSS.n17262 VSS.n14503 4.65
R14437 VSS.n17416 VSS.n17415 4.65
R14438 VSS.n17357 VSS.n17356 4.65
R14439 VSS.n17345 VSS.n17344 4.65
R14440 VSS.n17333 VSS.n17332 4.65
R14441 VSS.n17321 VSS.n17320 4.65
R14442 VSS.n17304 VSS.n17300 4.65
R14443 VSS.n17297 VSS.n17296 4.65
R14444 VSS.n17285 VSS.n17284 4.65
R14445 VSS.n17273 VSS.n17272 4.65
R14446 VSS.n17430 VSS.n14491 4.65
R14447 VSS.n17584 VSS.n17583 4.65
R14448 VSS.n17525 VSS.n17524 4.65
R14449 VSS.n17513 VSS.n17512 4.65
R14450 VSS.n17501 VSS.n17500 4.65
R14451 VSS.n17489 VSS.n17488 4.65
R14452 VSS.n17472 VSS.n17468 4.65
R14453 VSS.n17465 VSS.n17464 4.65
R14454 VSS.n17453 VSS.n17452 4.65
R14455 VSS.n17441 VSS.n17440 4.65
R14456 VSS.n14284 VSS.n14283 4.65
R14457 VSS.n14227 VSS.n14226 4.65
R14458 VSS.n14215 VSS.n14214 4.65
R14459 VSS.n14203 VSS.n14202 4.65
R14460 VSS.n14191 VSS.n14190 4.65
R14461 VSS.n14179 VSS.n14178 4.65
R14462 VSS.n14167 VSS.n14166 4.65
R14463 VSS.n14155 VSS.n14154 4.65
R14464 VSS.n14143 VSS.n14142 4.65
R14465 VSS.n14299 VSS.n14298 4.65
R14466 VSS.n14464 VSS.n14463 4.65
R14467 VSS.n14407 VSS.n14406 4.65
R14468 VSS.n14395 VSS.n14394 4.65
R14469 VSS.n14383 VSS.n14382 4.65
R14470 VSS.n14371 VSS.n14370 4.65
R14471 VSS.n14359 VSS.n14358 4.65
R14472 VSS.n14347 VSS.n14346 4.65
R14473 VSS.n14335 VSS.n14334 4.65
R14474 VSS.n14323 VSS.n14322 4.65
R14475 VSS.n14479 VSS.n14478 4.65
R14476 VSS.n12635 VSS.n12634 4.65
R14477 VSS.n10708 VSS.n10707 4.65
R14478 VSS.n10722 VSS.n10721 4.65
R14479 VSS.n10736 VSS.n10735 4.65
R14480 VSS.n10750 VSS.n10749 4.65
R14481 VSS.n10764 VSS.n10763 4.65
R14482 VSS.n10783 VSS.n10782 4.65
R14483 VSS.n10786 VSS.n10648 4.65
R14484 VSS.n10800 VSS.n10799 4.65
R14485 VSS.n10814 VSS.n10813 4.65
R14486 VSS.n10828 VSS.n10827 4.65
R14487 VSS.n10842 VSS.n10841 4.65
R14488 VSS.n10859 VSS.n10858 4.65
R14489 VSS.n10964 VSS.n10963 4.65
R14490 VSS.n10978 VSS.n10977 4.65
R14491 VSS.n10992 VSS.n10991 4.65
R14492 VSS.n11006 VSS.n11005 4.65
R14493 VSS.n11020 VSS.n11019 4.65
R14494 VSS.n11039 VSS.n11038 4.65
R14495 VSS.n11042 VSS.n10642 4.65
R14496 VSS.n11056 VSS.n11055 4.65
R14497 VSS.n11070 VSS.n11069 4.65
R14498 VSS.n11084 VSS.n11083 4.65
R14499 VSS.n11098 VSS.n11097 4.65
R14500 VSS.n11115 VSS.n11114 4.65
R14501 VSS.n11208 VSS.n11207 4.65
R14502 VSS.n11222 VSS.n11221 4.65
R14503 VSS.n11236 VSS.n11235 4.65
R14504 VSS.n11250 VSS.n11249 4.65
R14505 VSS.n11264 VSS.n11263 4.65
R14506 VSS.n11283 VSS.n11282 4.65
R14507 VSS.n11286 VSS.n10636 4.65
R14508 VSS.n11300 VSS.n11299 4.65
R14509 VSS.n11314 VSS.n11313 4.65
R14510 VSS.n11328 VSS.n11327 4.65
R14511 VSS.n11342 VSS.n11341 4.65
R14512 VSS.n11359 VSS.n11358 4.65
R14513 VSS.n11452 VSS.n11451 4.65
R14514 VSS.n11466 VSS.n11465 4.65
R14515 VSS.n11480 VSS.n11479 4.65
R14516 VSS.n11494 VSS.n11493 4.65
R14517 VSS.n11508 VSS.n11507 4.65
R14518 VSS.n11527 VSS.n11526 4.65
R14519 VSS.n11530 VSS.n10630 4.65
R14520 VSS.n11544 VSS.n11543 4.65
R14521 VSS.n11558 VSS.n11557 4.65
R14522 VSS.n11572 VSS.n11571 4.65
R14523 VSS.n11586 VSS.n11585 4.65
R14524 VSS.n11603 VSS.n11602 4.65
R14525 VSS.n11696 VSS.n11695 4.65
R14526 VSS.n11710 VSS.n11709 4.65
R14527 VSS.n11724 VSS.n11723 4.65
R14528 VSS.n11738 VSS.n11737 4.65
R14529 VSS.n11752 VSS.n11751 4.65
R14530 VSS.n11771 VSS.n11770 4.65
R14531 VSS.n11774 VSS.n10624 4.65
R14532 VSS.n11788 VSS.n11787 4.65
R14533 VSS.n11802 VSS.n11801 4.65
R14534 VSS.n11816 VSS.n11815 4.65
R14535 VSS.n11830 VSS.n11829 4.65
R14536 VSS.n11847 VSS.n11846 4.65
R14537 VSS.n11940 VSS.n11939 4.65
R14538 VSS.n11954 VSS.n11953 4.65
R14539 VSS.n11968 VSS.n11967 4.65
R14540 VSS.n11982 VSS.n11981 4.65
R14541 VSS.n11996 VSS.n11995 4.65
R14542 VSS.n12015 VSS.n12014 4.65
R14543 VSS.n12018 VSS.n10618 4.65
R14544 VSS.n12032 VSS.n12031 4.65
R14545 VSS.n12046 VSS.n12045 4.65
R14546 VSS.n12060 VSS.n12059 4.65
R14547 VSS.n12074 VSS.n12073 4.65
R14548 VSS.n12091 VSS.n12090 4.65
R14549 VSS.n12184 VSS.n12183 4.65
R14550 VSS.n12198 VSS.n12197 4.65
R14551 VSS.n12212 VSS.n12211 4.65
R14552 VSS.n12226 VSS.n12225 4.65
R14553 VSS.n12240 VSS.n12239 4.65
R14554 VSS.n12259 VSS.n12258 4.65
R14555 VSS.n12262 VSS.n10612 4.65
R14556 VSS.n12276 VSS.n12275 4.65
R14557 VSS.n12290 VSS.n12289 4.65
R14558 VSS.n12304 VSS.n12303 4.65
R14559 VSS.n12318 VSS.n12317 4.65
R14560 VSS.n12335 VSS.n12334 4.65
R14561 VSS.n12574 VSS.n12573 4.65
R14562 VSS.n12560 VSS.n12559 4.65
R14563 VSS.n12546 VSS.n12545 4.65
R14564 VSS.n12532 VSS.n12531 4.65
R14565 VSS.n12518 VSS.n10606 4.65
R14566 VSS.n12515 VSS.n12514 4.65
R14567 VSS.n12496 VSS.n12495 4.65
R14568 VSS.n12482 VSS.n12481 4.65
R14569 VSS.n12468 VSS.n12467 4.65
R14570 VSS.n12454 VSS.n12453 4.65
R14571 VSS.n12440 VSS.n12439 4.65
R14572 VSS.n12801 VSS.n12800 4.65
R14573 VSS.n12744 VSS.n12743 4.65
R14574 VSS.n12732 VSS.n12731 4.65
R14575 VSS.n12720 VSS.n12719 4.65
R14576 VSS.n12708 VSS.n12707 4.65
R14577 VSS.n12696 VSS.n12695 4.65
R14578 VSS.n12684 VSS.n12683 4.65
R14579 VSS.n12672 VSS.n12671 4.65
R14580 VSS.n12660 VSS.n12659 4.65
R14581 VSS.n12816 VSS.n12815 4.65
R14582 VSS.n12981 VSS.n12980 4.65
R14583 VSS.n12924 VSS.n12923 4.65
R14584 VSS.n12912 VSS.n12911 4.65
R14585 VSS.n12900 VSS.n12899 4.65
R14586 VSS.n12888 VSS.n12887 4.65
R14587 VSS.n12876 VSS.n12875 4.65
R14588 VSS.n12864 VSS.n12863 4.65
R14589 VSS.n12852 VSS.n12851 4.65
R14590 VSS.n12840 VSS.n12839 4.65
R14591 VSS.n12996 VSS.n12995 4.65
R14592 VSS.n13161 VSS.n13160 4.65
R14593 VSS.n13104 VSS.n13103 4.65
R14594 VSS.n13092 VSS.n13091 4.65
R14595 VSS.n13080 VSS.n13079 4.65
R14596 VSS.n13068 VSS.n13067 4.65
R14597 VSS.n13056 VSS.n13055 4.65
R14598 VSS.n13044 VSS.n13043 4.65
R14599 VSS.n13032 VSS.n13031 4.65
R14600 VSS.n13020 VSS.n13019 4.65
R14601 VSS.n13176 VSS.n13175 4.65
R14602 VSS.n13341 VSS.n13340 4.65
R14603 VSS.n13284 VSS.n13283 4.65
R14604 VSS.n13272 VSS.n13271 4.65
R14605 VSS.n13260 VSS.n13259 4.65
R14606 VSS.n13248 VSS.n13247 4.65
R14607 VSS.n13236 VSS.n13235 4.65
R14608 VSS.n13224 VSS.n13223 4.65
R14609 VSS.n13212 VSS.n13211 4.65
R14610 VSS.n13200 VSS.n13199 4.65
R14611 VSS.n13356 VSS.n13355 4.65
R14612 VSS.n13521 VSS.n13520 4.65
R14613 VSS.n13464 VSS.n13463 4.65
R14614 VSS.n13452 VSS.n13451 4.65
R14615 VSS.n13440 VSS.n13439 4.65
R14616 VSS.n13428 VSS.n13427 4.65
R14617 VSS.n13416 VSS.n13415 4.65
R14618 VSS.n13404 VSS.n13403 4.65
R14619 VSS.n13392 VSS.n13391 4.65
R14620 VSS.n13380 VSS.n13379 4.65
R14621 VSS.n13536 VSS.n13535 4.65
R14622 VSS.n13701 VSS.n13700 4.65
R14623 VSS.n13644 VSS.n13643 4.65
R14624 VSS.n13632 VSS.n13631 4.65
R14625 VSS.n13620 VSS.n13619 4.65
R14626 VSS.n13608 VSS.n13607 4.65
R14627 VSS.n13596 VSS.n13595 4.65
R14628 VSS.n13584 VSS.n13583 4.65
R14629 VSS.n13572 VSS.n13571 4.65
R14630 VSS.n13560 VSS.n13559 4.65
R14631 VSS.n13716 VSS.n13715 4.65
R14632 VSS.n13881 VSS.n13880 4.65
R14633 VSS.n13824 VSS.n13823 4.65
R14634 VSS.n13812 VSS.n13811 4.65
R14635 VSS.n13800 VSS.n13799 4.65
R14636 VSS.n13788 VSS.n13787 4.65
R14637 VSS.n13776 VSS.n13775 4.65
R14638 VSS.n13764 VSS.n13763 4.65
R14639 VSS.n13752 VSS.n13751 4.65
R14640 VSS.n13740 VSS.n13739 4.65
R14641 VSS.n13896 VSS.n13895 4.65
R14642 VSS.n14061 VSS.n14060 4.65
R14643 VSS.n14004 VSS.n14003 4.65
R14644 VSS.n13992 VSS.n13991 4.65
R14645 VSS.n13980 VSS.n13979 4.65
R14646 VSS.n13968 VSS.n13967 4.65
R14647 VSS.n13956 VSS.n13955 4.65
R14648 VSS.n13944 VSS.n13943 4.65
R14649 VSS.n13932 VSS.n13931 4.65
R14650 VSS.n13920 VSS.n13919 4.65
R14651 VSS.n9203 VSS.n9202 4.65
R14652 VSS.n7276 VSS.n7275 4.65
R14653 VSS.n7290 VSS.n7289 4.65
R14654 VSS.n7304 VSS.n7303 4.65
R14655 VSS.n7318 VSS.n7317 4.65
R14656 VSS.n7332 VSS.n7331 4.65
R14657 VSS.n7351 VSS.n7350 4.65
R14658 VSS.n7354 VSS.n7216 4.65
R14659 VSS.n7368 VSS.n7367 4.65
R14660 VSS.n7382 VSS.n7381 4.65
R14661 VSS.n7396 VSS.n7395 4.65
R14662 VSS.n7410 VSS.n7409 4.65
R14663 VSS.n7427 VSS.n7426 4.65
R14664 VSS.n7532 VSS.n7531 4.65
R14665 VSS.n7546 VSS.n7545 4.65
R14666 VSS.n7560 VSS.n7559 4.65
R14667 VSS.n7574 VSS.n7573 4.65
R14668 VSS.n7588 VSS.n7587 4.65
R14669 VSS.n7607 VSS.n7606 4.65
R14670 VSS.n7610 VSS.n7210 4.65
R14671 VSS.n7624 VSS.n7623 4.65
R14672 VSS.n7638 VSS.n7637 4.65
R14673 VSS.n7652 VSS.n7651 4.65
R14674 VSS.n7666 VSS.n7665 4.65
R14675 VSS.n7683 VSS.n7682 4.65
R14676 VSS.n7776 VSS.n7775 4.65
R14677 VSS.n7790 VSS.n7789 4.65
R14678 VSS.n7804 VSS.n7803 4.65
R14679 VSS.n7818 VSS.n7817 4.65
R14680 VSS.n7832 VSS.n7831 4.65
R14681 VSS.n7851 VSS.n7850 4.65
R14682 VSS.n7854 VSS.n7204 4.65
R14683 VSS.n7868 VSS.n7867 4.65
R14684 VSS.n7882 VSS.n7881 4.65
R14685 VSS.n7896 VSS.n7895 4.65
R14686 VSS.n7910 VSS.n7909 4.65
R14687 VSS.n7927 VSS.n7926 4.65
R14688 VSS.n8020 VSS.n8019 4.65
R14689 VSS.n8034 VSS.n8033 4.65
R14690 VSS.n8048 VSS.n8047 4.65
R14691 VSS.n8062 VSS.n8061 4.65
R14692 VSS.n8076 VSS.n8075 4.65
R14693 VSS.n8095 VSS.n8094 4.65
R14694 VSS.n8098 VSS.n7198 4.65
R14695 VSS.n8112 VSS.n8111 4.65
R14696 VSS.n8126 VSS.n8125 4.65
R14697 VSS.n8140 VSS.n8139 4.65
R14698 VSS.n8154 VSS.n8153 4.65
R14699 VSS.n8171 VSS.n8170 4.65
R14700 VSS.n8264 VSS.n8263 4.65
R14701 VSS.n8278 VSS.n8277 4.65
R14702 VSS.n8292 VSS.n8291 4.65
R14703 VSS.n8306 VSS.n8305 4.65
R14704 VSS.n8320 VSS.n8319 4.65
R14705 VSS.n8339 VSS.n8338 4.65
R14706 VSS.n8342 VSS.n7192 4.65
R14707 VSS.n8356 VSS.n8355 4.65
R14708 VSS.n8370 VSS.n8369 4.65
R14709 VSS.n8384 VSS.n8383 4.65
R14710 VSS.n8398 VSS.n8397 4.65
R14711 VSS.n8415 VSS.n8414 4.65
R14712 VSS.n8508 VSS.n8507 4.65
R14713 VSS.n8522 VSS.n8521 4.65
R14714 VSS.n8536 VSS.n8535 4.65
R14715 VSS.n8550 VSS.n8549 4.65
R14716 VSS.n8564 VSS.n8563 4.65
R14717 VSS.n8583 VSS.n8582 4.65
R14718 VSS.n8586 VSS.n7186 4.65
R14719 VSS.n8600 VSS.n8599 4.65
R14720 VSS.n8614 VSS.n8613 4.65
R14721 VSS.n8628 VSS.n8627 4.65
R14722 VSS.n8642 VSS.n8641 4.65
R14723 VSS.n8659 VSS.n8658 4.65
R14724 VSS.n8752 VSS.n8751 4.65
R14725 VSS.n8766 VSS.n8765 4.65
R14726 VSS.n8780 VSS.n8779 4.65
R14727 VSS.n8794 VSS.n8793 4.65
R14728 VSS.n8808 VSS.n8807 4.65
R14729 VSS.n8827 VSS.n8826 4.65
R14730 VSS.n8830 VSS.n7180 4.65
R14731 VSS.n8844 VSS.n8843 4.65
R14732 VSS.n8858 VSS.n8857 4.65
R14733 VSS.n8872 VSS.n8871 4.65
R14734 VSS.n8886 VSS.n8885 4.65
R14735 VSS.n8903 VSS.n8902 4.65
R14736 VSS.n9142 VSS.n9141 4.65
R14737 VSS.n9128 VSS.n9127 4.65
R14738 VSS.n9114 VSS.n9113 4.65
R14739 VSS.n9100 VSS.n9099 4.65
R14740 VSS.n9086 VSS.n7174 4.65
R14741 VSS.n9083 VSS.n9082 4.65
R14742 VSS.n9064 VSS.n9063 4.65
R14743 VSS.n9050 VSS.n9049 4.65
R14744 VSS.n9036 VSS.n9035 4.65
R14745 VSS.n9022 VSS.n9021 4.65
R14746 VSS.n9008 VSS.n9007 4.65
R14747 VSS.n10239 VSS.n10238 4.65
R14748 VSS.n10251 VSS.n10250 4.65
R14749 VSS.n10263 VSS.n10262 4.65
R14750 VSS.n10270 VSS.n10266 4.65
R14751 VSS.n10287 VSS.n10286 4.65
R14752 VSS.n10299 VSS.n10298 4.65
R14753 VSS.n10311 VSS.n10310 4.65
R14754 VSS.n10323 VSS.n10322 4.65
R14755 VSS.n10380 VSS.n10379 4.65
R14756 VSS.n10228 VSS.n10227 4.65
R14757 VSS.n10071 VSS.n10070 4.65
R14758 VSS.n10083 VSS.n10082 4.65
R14759 VSS.n10095 VSS.n10094 4.65
R14760 VSS.n10102 VSS.n10098 4.65
R14761 VSS.n10119 VSS.n10118 4.65
R14762 VSS.n10131 VSS.n10130 4.65
R14763 VSS.n10143 VSS.n10142 4.65
R14764 VSS.n10155 VSS.n10154 4.65
R14765 VSS.n10212 VSS.n10211 4.65
R14766 VSS.n10060 VSS.n10059 4.65
R14767 VSS.n9903 VSS.n9902 4.65
R14768 VSS.n9915 VSS.n9914 4.65
R14769 VSS.n9927 VSS.n9926 4.65
R14770 VSS.n9934 VSS.n9930 4.65
R14771 VSS.n9951 VSS.n9950 4.65
R14772 VSS.n9963 VSS.n9962 4.65
R14773 VSS.n9975 VSS.n9974 4.65
R14774 VSS.n9987 VSS.n9986 4.65
R14775 VSS.n10044 VSS.n10043 4.65
R14776 VSS.n9892 VSS.n9891 4.65
R14777 VSS.n9735 VSS.n9734 4.65
R14778 VSS.n9747 VSS.n9746 4.65
R14779 VSS.n9759 VSS.n9758 4.65
R14780 VSS.n9766 VSS.n9762 4.65
R14781 VSS.n9783 VSS.n9782 4.65
R14782 VSS.n9795 VSS.n9794 4.65
R14783 VSS.n9807 VSS.n9806 4.65
R14784 VSS.n9819 VSS.n9818 4.65
R14785 VSS.n9876 VSS.n9875 4.65
R14786 VSS.n9724 VSS.n9723 4.65
R14787 VSS.n9567 VSS.n9566 4.65
R14788 VSS.n9579 VSS.n9578 4.65
R14789 VSS.n9591 VSS.n9590 4.65
R14790 VSS.n9598 VSS.n9594 4.65
R14791 VSS.n9615 VSS.n9614 4.65
R14792 VSS.n9627 VSS.n9626 4.65
R14793 VSS.n9639 VSS.n9638 4.65
R14794 VSS.n9651 VSS.n9650 4.65
R14795 VSS.n9708 VSS.n9707 4.65
R14796 VSS.n9556 VSS.n9555 4.65
R14797 VSS.n9399 VSS.n9398 4.65
R14798 VSS.n9411 VSS.n9410 4.65
R14799 VSS.n9423 VSS.n9422 4.65
R14800 VSS.n9430 VSS.n9426 4.65
R14801 VSS.n9447 VSS.n9446 4.65
R14802 VSS.n9459 VSS.n9458 4.65
R14803 VSS.n9471 VSS.n9470 4.65
R14804 VSS.n9483 VSS.n9482 4.65
R14805 VSS.n9540 VSS.n9539 4.65
R14806 VSS.n9388 VSS.n9387 4.65
R14807 VSS.n9231 VSS.n9230 4.65
R14808 VSS.n9243 VSS.n9242 4.65
R14809 VSS.n9255 VSS.n9254 4.65
R14810 VSS.n9262 VSS.n9258 4.65
R14811 VSS.n9279 VSS.n9278 4.65
R14812 VSS.n9291 VSS.n9290 4.65
R14813 VSS.n9303 VSS.n9302 4.65
R14814 VSS.n9315 VSS.n9314 4.65
R14815 VSS.n9372 VSS.n9371 4.65
R14816 VSS.n9220 VSS.n9219 4.65
R14817 VSS.n10548 VSS.n10547 4.65
R14818 VSS.n10490 VSS.n10489 4.65
R14819 VSS.n10478 VSS.n10477 4.65
R14820 VSS.n10466 VSS.n10465 4.65
R14821 VSS.n10454 VSS.n10453 4.65
R14822 VSS.n10437 VSS.n10433 4.65
R14823 VSS.n10430 VSS.n10429 4.65
R14824 VSS.n10418 VSS.n10417 4.65
R14825 VSS.n10406 VSS.n10405 4.65
R14826 VSS.n10395 VSS.n10394 4.65
R14827 VSS.n4838 VSS.n4837 4.65
R14828 VSS.n3459 VSS.n3452 4.65
R14829 VSS.n3797 VSS.n3458 4.65
R14830 VSS.n3787 VSS.n3786 4.65
R14831 VSS.n3471 VSS.n3468 4.65
R14832 VSS.n3774 VSS.n3478 4.65
R14833 VSS.n3764 VSS.n3763 4.65
R14834 VSS.n3490 VSS.n3487 4.65
R14835 VSS.n3751 VSS.n3497 4.65
R14836 VSS.n3741 VSS.n3740 4.65
R14837 VSS.n3509 VSS.n3506 4.65
R14838 VSS.n3728 VSS.n3516 4.65
R14839 VSS.n3718 VSS.n3717 4.65
R14840 VSS.n3561 VSS.n3559 4.65
R14841 VSS.n3704 VSS.n3571 4.65
R14842 VSS.n3694 VSS.n3693 4.65
R14843 VSS.n3583 VSS.n3580 4.65
R14844 VSS.n3681 VSS.n3590 4.65
R14845 VSS.n3671 VSS.n3670 4.65
R14846 VSS.n3602 VSS.n3599 4.65
R14847 VSS.n3658 VSS.n3609 4.65
R14848 VSS.n3648 VSS.n3647 4.65
R14849 VSS.n3621 VSS.n3618 4.65
R14850 VSS.n3635 VSS.n3632 4.65
R14851 VSS.n3954 VSS.n3390 4.65
R14852 VSS.n3966 VSS.n3381 4.65
R14853 VSS.n3976 VSS.n3375 4.65
R14854 VSS.n3370 VSS.n3369 4.65
R14855 VSS.n3990 VSS.n3368 4.65
R14856 VSS.n4001 VSS.n3360 4.65
R14857 VSS.n4011 VSS.n3354 4.65
R14858 VSS.n3349 VSS.n3348 4.65
R14859 VSS.n4025 VSS.n3347 4.65
R14860 VSS.n4036 VSS.n3339 4.65
R14861 VSS.n4046 VSS.n3333 4.65
R14862 VSS.n3328 VSS.n3327 4.65
R14863 VSS.n4415 VSS.n3326 4.65
R14864 VSS.n4062 VSS.n4060 4.65
R14865 VSS.n4401 VSS.n4071 4.65
R14866 VSS.n4391 VSS.n4390 4.65
R14867 VSS.n4083 VSS.n4080 4.65
R14868 VSS.n4378 VSS.n4090 4.65
R14869 VSS.n4368 VSS.n4367 4.65
R14870 VSS.n4102 VSS.n4099 4.65
R14871 VSS.n4355 VSS.n4109 4.65
R14872 VSS.n4345 VSS.n4344 4.65
R14873 VSS.n4121 VSS.n4118 4.65
R14874 VSS.n4332 VSS.n4128 4.65
R14875 VSS.n4322 VSS.n4321 4.65
R14876 VSS.n4173 VSS.n4171 4.65
R14877 VSS.n4308 VSS.n4183 4.65
R14878 VSS.n4298 VSS.n4297 4.65
R14879 VSS.n4195 VSS.n4192 4.65
R14880 VSS.n4285 VSS.n4202 4.65
R14881 VSS.n4275 VSS.n4274 4.65
R14882 VSS.n4214 VSS.n4211 4.65
R14883 VSS.n4262 VSS.n4221 4.65
R14884 VSS.n4252 VSS.n4251 4.65
R14885 VSS.n4233 VSS.n4230 4.65
R14886 VSS.n3223 VSS.n3222 4.65
R14887 VSS.n4541 VSS.n4540 4.65
R14888 VSS.n3214 VSS.n3213 4.65
R14889 VSS.n4556 VSS.n3212 4.65
R14890 VSS.n4567 VSS.n3204 4.65
R14891 VSS.n4577 VSS.n3198 4.65
R14892 VSS.n3193 VSS.n3192 4.65
R14893 VSS.n4591 VSS.n3191 4.65
R14894 VSS.n4602 VSS.n3183 4.65
R14895 VSS.n4612 VSS.n3177 4.65
R14896 VSS.n3172 VSS.n3171 4.65
R14897 VSS.n4626 VSS.n3170 4.65
R14898 VSS.n4637 VSS.n3162 4.65
R14899 VSS.n4648 VSS.n4647 4.65
R14900 VSS.n4652 VSS.n4650 4.65
R14901 VSS.n5010 VSS.n4661 4.65
R14902 VSS.n5000 VSS.n4999 4.65
R14903 VSS.n4673 VSS.n4670 4.65
R14904 VSS.n4987 VSS.n4680 4.65
R14905 VSS.n4977 VSS.n4976 4.65
R14906 VSS.n4692 VSS.n4689 4.65
R14907 VSS.n4964 VSS.n4699 4.65
R14908 VSS.n4954 VSS.n4953 4.65
R14909 VSS.n4711 VSS.n4708 4.65
R14910 VSS.n4941 VSS.n4718 4.65
R14911 VSS.n4931 VSS.n4930 4.65
R14912 VSS.n4848 VSS.n4830 4.65
R14913 VSS.n4823 VSS.n4820 4.65
R14914 VSS.n4861 VSS.n4860 4.65
R14915 VSS.n4871 VSS.n4811 4.65
R14916 VSS.n4804 VSS.n4801 4.65
R14917 VSS.n4884 VSS.n4883 4.65
R14918 VSS.n4894 VSS.n4792 4.65
R14919 VSS.n4785 VSS.n4782 4.65
R14920 VSS.n4907 VSS.n4906 4.65
R14921 VSS.n4917 VSS.n4773 4.65
R14922 VSS.n4763 VSS.n4761 4.65
R14923 VSS.n3038 VSS.n3034 4.65
R14924 VSS.n3049 VSS.n3028 4.65
R14925 VSS.n3054 VSS.n3025 4.65
R14926 VSS.n3060 VSS.n3021 4.65
R14927 VSS.n3066 VSS.n3015 4.65
R14928 VSS.n3072 VSS.n3071 4.65
R14929 VSS.n3080 VSS.n1695 4.65
R14930 VSS.n2948 VSS.n2944 4.65
R14931 VSS.n2959 VSS.n2938 4.65
R14932 VSS.n2964 VSS.n2935 4.65
R14933 VSS.n2970 VSS.n2931 4.65
R14934 VSS.n2976 VSS.n2925 4.65
R14935 VSS.n2982 VSS.n2981 4.65
R14936 VSS.n2990 VSS.n1785 4.65
R14937 VSS.n2858 VSS.n2854 4.65
R14938 VSS.n2869 VSS.n2848 4.65
R14939 VSS.n2874 VSS.n2845 4.65
R14940 VSS.n2880 VSS.n2841 4.65
R14941 VSS.n2886 VSS.n2835 4.65
R14942 VSS.n2892 VSS.n2891 4.65
R14943 VSS.n2900 VSS.n1875 4.65
R14944 VSS.n2768 VSS.n2764 4.65
R14945 VSS.n2779 VSS.n2758 4.65
R14946 VSS.n2784 VSS.n2755 4.65
R14947 VSS.n2790 VSS.n2751 4.65
R14948 VSS.n2796 VSS.n2745 4.65
R14949 VSS.n2802 VSS.n2801 4.65
R14950 VSS.n2810 VSS.n1965 4.65
R14951 VSS.n2678 VSS.n2674 4.65
R14952 VSS.n2689 VSS.n2668 4.65
R14953 VSS.n2694 VSS.n2665 4.65
R14954 VSS.n2700 VSS.n2661 4.65
R14955 VSS.n2706 VSS.n2655 4.65
R14956 VSS.n2712 VSS.n2711 4.65
R14957 VSS.n2720 VSS.n2055 4.65
R14958 VSS.n2588 VSS.n2584 4.65
R14959 VSS.n2599 VSS.n2578 4.65
R14960 VSS.n2604 VSS.n2575 4.65
R14961 VSS.n2610 VSS.n2571 4.65
R14962 VSS.n2616 VSS.n2565 4.65
R14963 VSS.n2622 VSS.n2621 4.65
R14964 VSS.n2630 VSS.n2145 4.65
R14965 VSS.n2498 VSS.n2494 4.65
R14966 VSS.n2509 VSS.n2488 4.65
R14967 VSS.n2514 VSS.n2485 4.65
R14968 VSS.n2520 VSS.n2481 4.65
R14969 VSS.n2526 VSS.n2475 4.65
R14970 VSS.n2532 VSS.n2531 4.65
R14971 VSS.n2540 VSS.n2235 4.65
R14972 VSS.n2408 VSS.n2404 4.65
R14973 VSS.n2419 VSS.n2398 4.65
R14974 VSS.n2424 VSS.n2395 4.65
R14975 VSS.n2430 VSS.n2391 4.65
R14976 VSS.n2436 VSS.n2385 4.65
R14977 VSS.n2442 VSS.n2441 4.65
R14978 VSS.n2450 VSS.n2325 4.65
R14979 VSS.n2381 VSS.n2380 4.65
R14980 VSS.n2413 VSS.n2401 4.65
R14981 VSS.n2463 VSS.n2462 4.65
R14982 VSS.n2471 VSS.n2470 4.65
R14983 VSS.n2503 VSS.n2491 4.65
R14984 VSS.n2553 VSS.n2552 4.65
R14985 VSS.n2561 VSS.n2560 4.65
R14986 VSS.n2593 VSS.n2581 4.65
R14987 VSS.n2643 VSS.n2642 4.65
R14988 VSS.n2651 VSS.n2650 4.65
R14989 VSS.n2683 VSS.n2671 4.65
R14990 VSS.n2733 VSS.n2732 4.65
R14991 VSS.n2741 VSS.n2740 4.65
R14992 VSS.n2773 VSS.n2761 4.65
R14993 VSS.n2823 VSS.n2822 4.65
R14994 VSS.n2831 VSS.n2830 4.65
R14995 VSS.n2863 VSS.n2851 4.65
R14996 VSS.n2913 VSS.n2912 4.65
R14997 VSS.n2921 VSS.n2920 4.65
R14998 VSS.n2953 VSS.n2941 4.65
R14999 VSS.n3003 VSS.n3002 4.65
R15000 VSS.n3011 VSS.n3010 4.65
R15001 VSS.n3043 VSS.n3031 4.65
R15002 VSS.n3093 VSS.n3092 4.65
R15003 VSS.n5134 VSS.n5133 4.65
R15004 VSS.n1171 VSS.n1170 4.65
R15005 VSS.n5142 VSS.n1581 4.65
R15006 VSS.n1576 VSS.n1575 4.65
R15007 VSS.n5156 VSS.n1574 4.65
R15008 VSS.n5167 VSS.n1566 4.65
R15009 VSS.n5177 VSS.n1560 4.65
R15010 VSS.n1555 VSS.n1554 4.65
R15011 VSS.n5191 VSS.n1553 4.65
R15012 VSS.n5202 VSS.n1545 4.65
R15013 VSS.n5212 VSS.n1539 4.65
R15014 VSS.n1532 VSS.n1531 4.65
R15015 VSS.n5229 VSS.n5228 4.65
R15016 VSS.n5406 VSS.n1523 4.65
R15017 VSS.n5394 VSS.n5237 4.65
R15018 VSS.n5384 VSS.n5383 4.65
R15019 VSS.n5248 VSS.n5245 4.65
R15020 VSS.n5371 VSS.n5255 4.65
R15021 VSS.n5361 VSS.n5360 4.65
R15022 VSS.n5267 VSS.n5264 4.65
R15023 VSS.n5348 VSS.n5274 4.65
R15024 VSS.n5338 VSS.n5337 4.65
R15025 VSS.n5286 VSS.n5283 4.65
R15026 VSS.n5325 VSS.n5293 4.65
R15027 VSS.n5315 VSS.n5314 4.65
R15028 VSS.n5306 VSS.n5303 4.65
R15029 VSS.n5501 VSS.n1440 4.65
R15030 VSS.n1435 VSS.n1434 4.65
R15031 VSS.n5515 VSS.n1433 4.65
R15032 VSS.n5526 VSS.n1425 4.65
R15033 VSS.n5536 VSS.n1419 4.65
R15034 VSS.n1414 VSS.n1413 4.65
R15035 VSS.n5550 VSS.n1412 4.65
R15036 VSS.n5561 VSS.n1404 4.65
R15037 VSS.n5571 VSS.n1398 4.65
R15038 VSS.n1391 VSS.n1390 4.65
R15039 VSS.n5588 VSS.n5587 4.65
R15040 VSS.n5614 VSS.n1382 4.65
R15041 VSS.n5602 VSS.n5601 4.65
R15042 VSS.n522 VSS.n520 4.65
R15043 VSS.n5773 VSS.n529 4.65
R15044 VSS.n5763 VSS.n5762 4.65
R15045 VSS.n541 VSS.n538 4.65
R15046 VSS.n5750 VSS.n548 4.65
R15047 VSS.n5740 VSS.n5739 4.65
R15048 VSS.n560 VSS.n557 4.65
R15049 VSS.n5727 VSS.n567 4.65
R15050 VSS.n5717 VSS.n5716 4.65
R15051 VSS.n579 VSS.n576 4.65
R15052 VSS.n5704 VSS.n586 4.65
R15053 VSS.n787 VSS.n777 4.65
R15054 VSS.n772 VSS.n771 4.65
R15055 VSS.n801 VSS.n770 4.65
R15056 VSS.n812 VSS.n762 4.65
R15057 VSS.n822 VSS.n756 4.65
R15058 VSS.n751 VSS.n750 4.65
R15059 VSS.n836 VSS.n749 4.65
R15060 VSS.n847 VSS.n741 4.65
R15061 VSS.n857 VSS.n735 4.65
R15062 VSS.n730 VSS.n729 4.65
R15063 VSS.n871 VSS.n728 4.65
R15064 VSS.n882 VSS.n719 4.65
R15065 VSS.n924 VSS.n711 4.65
R15066 VSS.n934 VSS.n705 4.65
R15067 VSS.n700 VSS.n699 4.65
R15068 VSS.n948 VSS.n698 4.65
R15069 VSS.n959 VSS.n690 4.65
R15070 VSS.n969 VSS.n684 4.65
R15071 VSS.n679 VSS.n678 4.65
R15072 VSS.n983 VSS.n677 4.65
R15073 VSS.n994 VSS.n669 4.65
R15074 VSS.n1004 VSS.n663 4.65
R15075 VSS.n658 VSS.n657 4.65
R15076 VSS.n1264 VSS.n656 4.65
R15077 VSS.n1181 VSS.n1086 4.65
R15078 VSS.n1079 VSS.n1076 4.65
R15079 VSS.n1194 VSS.n1193 4.65
R15080 VSS.n1204 VSS.n1067 4.65
R15081 VSS.n1060 VSS.n1057 4.65
R15082 VSS.n1217 VSS.n1216 4.65
R15083 VSS.n1227 VSS.n1048 4.65
R15084 VSS.n1041 VSS.n1038 4.65
R15085 VSS.n1240 VSS.n1239 4.65
R15086 VSS.n1250 VSS.n1029 4.65
R15087 VSS.n1020 VSS.n1018 4.65
R15088 VSS.n6701 VSS.n6699 4.65
R15089 VSS.n6706 VSS.n6696 4.65
R15090 VSS.n6711 VSS.n6693 4.65
R15091 VSS.n6717 VSS.n6689 4.65
R15092 VSS.n6723 VSS.n6685 4.65
R15093 VSS.n6729 VSS.n6679 4.65
R15094 VSS.n6735 VSS.n6734 4.65
R15095 VSS.n6743 VSS.n6619 4.65
R15096 VSS.n6675 VSS.n6674 4.65
R15097 VSS.n6757 VSS.n6756 4.65
R15098 VSS.n6791 VSS.n6789 4.65
R15099 VSS.n6796 VSS.n6786 4.65
R15100 VSS.n6801 VSS.n6783 4.65
R15101 VSS.n6807 VSS.n6779 4.65
R15102 VSS.n6813 VSS.n6775 4.65
R15103 VSS.n6819 VSS.n6769 4.65
R15104 VSS.n6825 VSS.n6824 4.65
R15105 VSS.n6833 VSS.n6529 4.65
R15106 VSS.n6765 VSS.n6764 4.65
R15107 VSS.n6847 VSS.n6846 4.65
R15108 VSS.n6881 VSS.n6879 4.65
R15109 VSS.n6886 VSS.n6876 4.65
R15110 VSS.n6891 VSS.n6873 4.65
R15111 VSS.n6897 VSS.n6869 4.65
R15112 VSS.n6903 VSS.n6865 4.65
R15113 VSS.n6909 VSS.n6859 4.65
R15114 VSS.n6915 VSS.n6914 4.65
R15115 VSS.n6923 VSS.n6439 4.65
R15116 VSS.n6855 VSS.n6854 4.65
R15117 VSS.n6937 VSS.n6936 4.65
R15118 VSS.n6128 VSS.n6125 4.65
R15119 VSS.n6136 VSS.n6123 4.65
R15120 VSS.n6144 VSS.n6121 4.65
R15121 VSS.n6152 VSS.n6119 4.65
R15122 VSS.n6160 VSS.n6117 4.65
R15123 VSS.n6168 VSS.n6115 4.65
R15124 VSS.n6176 VSS.n6113 4.65
R15125 VSS.n6184 VSS.n6111 4.65
R15126 VSS.n6243 VSS.n6110 4.65
R15127 VSS.n6240 VSS.n6189 4.65
R15128 VSS.n6012 VSS.n6009 4.65
R15129 VSS.n6020 VSS.n6007 4.65
R15130 VSS.n6028 VSS.n6005 4.65
R15131 VSS.n6036 VSS.n6003 4.65
R15132 VSS.n6044 VSS.n6001 4.65
R15133 VSS.n6052 VSS.n5999 4.65
R15134 VSS.n6060 VSS.n5997 4.65
R15135 VSS.n6068 VSS.n5995 4.65
R15136 VSS.n6307 VSS.n5994 4.65
R15137 VSS.n6304 VSS.n6253 4.65
R15138 VSS.n5896 VSS.n5893 4.65
R15139 VSS.n5904 VSS.n5891 4.65
R15140 VSS.n5912 VSS.n5889 4.65
R15141 VSS.n5920 VSS.n5887 4.65
R15142 VSS.n5928 VSS.n5885 4.65
R15143 VSS.n5936 VSS.n5883 4.65
R15144 VSS.n5944 VSS.n5881 4.65
R15145 VSS.n5952 VSS.n5879 4.65
R15146 VSS.n6371 VSS.n5878 4.65
R15147 VSS.n6368 VSS.n6317 4.65
R15148 VSS.n5788 VSS.n5786 4.65
R15149 VSS.n5798 VSS.n5792 4.65
R15150 VSS.n5804 VSS.n5797 4.65
R15151 VSS.n5810 VSS.n5803 4.65
R15152 VSS.n5815 VSS.n5809 4.65
R15153 VSS.n5822 VSS.n5821 4.65
R15154 VSS.n5828 VSS.n5820 4.65
R15155 VSS.n5834 VSS.n5827 4.65
R15156 VSS.n5839 VSS.n5833 4.65
R15157 VSS.n6382 VSS.n6381 4.65
R15158 VSS.n409 VSS.n408 4.65
R15159 VSS.n18023 VSS.n17921 4.65
R15160 VSS.n18201 VSS.n18200 4.65
R15161 VSS.n16375 VSS.n16374 4.608
R15162 VSS.n16374 VSS.n16371 4.608
R15163 VSS.n16371 VSS.n16368 4.608
R15164 VSS.n16368 VSS.n16365 4.608
R15165 VSS.n16365 VSS.n16362 4.608
R15166 VSS.n16362 VSS.n16359 4.608
R15167 VSS.n16359 VSS.n16356 4.608
R15168 VSS.n16356 VSS.n16353 4.608
R15169 VSS.n16353 VSS.n16350 4.608
R15170 VSS.n16350 VSS.n16347 4.608
R15171 VSS.n16347 VSS.n16344 4.608
R15172 VSS.n16344 VSS.n16341 4.608
R15173 VSS.n16120 VSS.n16119 4.608
R15174 VSS.n16119 VSS.n16116 4.608
R15175 VSS.n16116 VSS.n16113 4.608
R15176 VSS.n16113 VSS.n16110 4.608
R15177 VSS.n16110 VSS.n16107 4.608
R15178 VSS.n16107 VSS.n16104 4.608
R15179 VSS.n16104 VSS.n16101 4.608
R15180 VSS.n16101 VSS.n16098 4.608
R15181 VSS.n16098 VSS.n16095 4.608
R15182 VSS.n16095 VSS.n16092 4.608
R15183 VSS.n16092 VSS.n16089 4.608
R15184 VSS.n16089 VSS.n16086 4.608
R15185 VSS.n15875 VSS.n15874 4.608
R15186 VSS.n15874 VSS.n15871 4.608
R15187 VSS.n15871 VSS.n15868 4.608
R15188 VSS.n15868 VSS.n15865 4.608
R15189 VSS.n15865 VSS.n15862 4.608
R15190 VSS.n15862 VSS.n15859 4.608
R15191 VSS.n15859 VSS.n15856 4.608
R15192 VSS.n15856 VSS.n15853 4.608
R15193 VSS.n15853 VSS.n15850 4.608
R15194 VSS.n15850 VSS.n15847 4.608
R15195 VSS.n15847 VSS.n15844 4.608
R15196 VSS.n15844 VSS.n15841 4.608
R15197 VSS.n15632 VSS.n15631 4.608
R15198 VSS.n15631 VSS.n15628 4.608
R15199 VSS.n15628 VSS.n15625 4.608
R15200 VSS.n15625 VSS.n15622 4.608
R15201 VSS.n15622 VSS.n15619 4.608
R15202 VSS.n15619 VSS.n15616 4.608
R15203 VSS.n15616 VSS.n15613 4.608
R15204 VSS.n15613 VSS.n15610 4.608
R15205 VSS.n15610 VSS.n15607 4.608
R15206 VSS.n15607 VSS.n15604 4.608
R15207 VSS.n15604 VSS.n15601 4.608
R15208 VSS.n15601 VSS.n15598 4.608
R15209 VSS.n15387 VSS.n15386 4.608
R15210 VSS.n15386 VSS.n15383 4.608
R15211 VSS.n15383 VSS.n15380 4.608
R15212 VSS.n15380 VSS.n15377 4.608
R15213 VSS.n15377 VSS.n15374 4.608
R15214 VSS.n15374 VSS.n15371 4.608
R15215 VSS.n15371 VSS.n15368 4.608
R15216 VSS.n15368 VSS.n15365 4.608
R15217 VSS.n15365 VSS.n15362 4.608
R15218 VSS.n15362 VSS.n15359 4.608
R15219 VSS.n15359 VSS.n15356 4.608
R15220 VSS.n15356 VSS.n15353 4.608
R15221 VSS.n15144 VSS.n15143 4.608
R15222 VSS.n15143 VSS.n15140 4.608
R15223 VSS.n15140 VSS.n15137 4.608
R15224 VSS.n15137 VSS.n15134 4.608
R15225 VSS.n15134 VSS.n15131 4.608
R15226 VSS.n15131 VSS.n15128 4.608
R15227 VSS.n15128 VSS.n15125 4.608
R15228 VSS.n15125 VSS.n15122 4.608
R15229 VSS.n15122 VSS.n15119 4.608
R15230 VSS.n15119 VSS.n15116 4.608
R15231 VSS.n15116 VSS.n15113 4.608
R15232 VSS.n15113 VSS.n15110 4.608
R15233 VSS.n14899 VSS.n14898 4.608
R15234 VSS.n14898 VSS.n14895 4.608
R15235 VSS.n14895 VSS.n14892 4.608
R15236 VSS.n14892 VSS.n14889 4.608
R15237 VSS.n14889 VSS.n14886 4.608
R15238 VSS.n14886 VSS.n14883 4.608
R15239 VSS.n14883 VSS.n14880 4.608
R15240 VSS.n14880 VSS.n14877 4.608
R15241 VSS.n14877 VSS.n14874 4.608
R15242 VSS.n14874 VSS.n14871 4.608
R15243 VSS.n14871 VSS.n14868 4.608
R15244 VSS.n14868 VSS.n14865 4.608
R15245 VSS.n12424 VSS.n12423 4.608
R15246 VSS.n12423 VSS.n12420 4.608
R15247 VSS.n12420 VSS.n12417 4.608
R15248 VSS.n12417 VSS.n12414 4.608
R15249 VSS.n12414 VSS.n12411 4.608
R15250 VSS.n12411 VSS.n12408 4.608
R15251 VSS.n12408 VSS.n12405 4.608
R15252 VSS.n12405 VSS.n12402 4.608
R15253 VSS.n12402 VSS.n12399 4.608
R15254 VSS.n12399 VSS.n12396 4.608
R15255 VSS.n12396 VSS.n12393 4.608
R15256 VSS.n12393 VSS.n12390 4.608
R15257 VSS.n12169 VSS.n12168 4.608
R15258 VSS.n12168 VSS.n12165 4.608
R15259 VSS.n12165 VSS.n12162 4.608
R15260 VSS.n12162 VSS.n12159 4.608
R15261 VSS.n12159 VSS.n12156 4.608
R15262 VSS.n12156 VSS.n12153 4.608
R15263 VSS.n12153 VSS.n12150 4.608
R15264 VSS.n12150 VSS.n12147 4.608
R15265 VSS.n12147 VSS.n12144 4.608
R15266 VSS.n12144 VSS.n12141 4.608
R15267 VSS.n12141 VSS.n12138 4.608
R15268 VSS.n12138 VSS.n12135 4.608
R15269 VSS.n11924 VSS.n11923 4.608
R15270 VSS.n11923 VSS.n11920 4.608
R15271 VSS.n11920 VSS.n11917 4.608
R15272 VSS.n11917 VSS.n11914 4.608
R15273 VSS.n11914 VSS.n11911 4.608
R15274 VSS.n11911 VSS.n11908 4.608
R15275 VSS.n11908 VSS.n11905 4.608
R15276 VSS.n11905 VSS.n11902 4.608
R15277 VSS.n11902 VSS.n11899 4.608
R15278 VSS.n11899 VSS.n11896 4.608
R15279 VSS.n11896 VSS.n11893 4.608
R15280 VSS.n11893 VSS.n11890 4.608
R15281 VSS.n11681 VSS.n11680 4.608
R15282 VSS.n11680 VSS.n11677 4.608
R15283 VSS.n11677 VSS.n11674 4.608
R15284 VSS.n11674 VSS.n11671 4.608
R15285 VSS.n11671 VSS.n11668 4.608
R15286 VSS.n11668 VSS.n11665 4.608
R15287 VSS.n11665 VSS.n11662 4.608
R15288 VSS.n11662 VSS.n11659 4.608
R15289 VSS.n11659 VSS.n11656 4.608
R15290 VSS.n11656 VSS.n11653 4.608
R15291 VSS.n11653 VSS.n11650 4.608
R15292 VSS.n11650 VSS.n11647 4.608
R15293 VSS.n11436 VSS.n11435 4.608
R15294 VSS.n11435 VSS.n11432 4.608
R15295 VSS.n11432 VSS.n11429 4.608
R15296 VSS.n11429 VSS.n11426 4.608
R15297 VSS.n11426 VSS.n11423 4.608
R15298 VSS.n11423 VSS.n11420 4.608
R15299 VSS.n11420 VSS.n11417 4.608
R15300 VSS.n11417 VSS.n11414 4.608
R15301 VSS.n11414 VSS.n11411 4.608
R15302 VSS.n11411 VSS.n11408 4.608
R15303 VSS.n11408 VSS.n11405 4.608
R15304 VSS.n11405 VSS.n11402 4.608
R15305 VSS.n11193 VSS.n11192 4.608
R15306 VSS.n11192 VSS.n11189 4.608
R15307 VSS.n11189 VSS.n11186 4.608
R15308 VSS.n11186 VSS.n11183 4.608
R15309 VSS.n11183 VSS.n11180 4.608
R15310 VSS.n11180 VSS.n11177 4.608
R15311 VSS.n11177 VSS.n11174 4.608
R15312 VSS.n11174 VSS.n11171 4.608
R15313 VSS.n11171 VSS.n11168 4.608
R15314 VSS.n11168 VSS.n11165 4.608
R15315 VSS.n11165 VSS.n11162 4.608
R15316 VSS.n11162 VSS.n11159 4.608
R15317 VSS.n10948 VSS.n10947 4.608
R15318 VSS.n10947 VSS.n10944 4.608
R15319 VSS.n10944 VSS.n10941 4.608
R15320 VSS.n10941 VSS.n10938 4.608
R15321 VSS.n10938 VSS.n10935 4.608
R15322 VSS.n10935 VSS.n10932 4.608
R15323 VSS.n10932 VSS.n10929 4.608
R15324 VSS.n10929 VSS.n10926 4.608
R15325 VSS.n10926 VSS.n10923 4.608
R15326 VSS.n10923 VSS.n10920 4.608
R15327 VSS.n10920 VSS.n10917 4.608
R15328 VSS.n10917 VSS.n10914 4.608
R15329 VSS.n8992 VSS.n8991 4.608
R15330 VSS.n8991 VSS.n8988 4.608
R15331 VSS.n8988 VSS.n8985 4.608
R15332 VSS.n8985 VSS.n8982 4.608
R15333 VSS.n8982 VSS.n8979 4.608
R15334 VSS.n8979 VSS.n8976 4.608
R15335 VSS.n8976 VSS.n8973 4.608
R15336 VSS.n8973 VSS.n8970 4.608
R15337 VSS.n8970 VSS.n8967 4.608
R15338 VSS.n8967 VSS.n8964 4.608
R15339 VSS.n8964 VSS.n8961 4.608
R15340 VSS.n8961 VSS.n8958 4.608
R15341 VSS.n8737 VSS.n8736 4.608
R15342 VSS.n8736 VSS.n8733 4.608
R15343 VSS.n8733 VSS.n8730 4.608
R15344 VSS.n8730 VSS.n8727 4.608
R15345 VSS.n8727 VSS.n8724 4.608
R15346 VSS.n8724 VSS.n8721 4.608
R15347 VSS.n8721 VSS.n8718 4.608
R15348 VSS.n8718 VSS.n8715 4.608
R15349 VSS.n8715 VSS.n8712 4.608
R15350 VSS.n8712 VSS.n8709 4.608
R15351 VSS.n8709 VSS.n8706 4.608
R15352 VSS.n8706 VSS.n8703 4.608
R15353 VSS.n8492 VSS.n8491 4.608
R15354 VSS.n8491 VSS.n8488 4.608
R15355 VSS.n8488 VSS.n8485 4.608
R15356 VSS.n8485 VSS.n8482 4.608
R15357 VSS.n8482 VSS.n8479 4.608
R15358 VSS.n8479 VSS.n8476 4.608
R15359 VSS.n8476 VSS.n8473 4.608
R15360 VSS.n8473 VSS.n8470 4.608
R15361 VSS.n8470 VSS.n8467 4.608
R15362 VSS.n8467 VSS.n8464 4.608
R15363 VSS.n8464 VSS.n8461 4.608
R15364 VSS.n8461 VSS.n8458 4.608
R15365 VSS.n8249 VSS.n8248 4.608
R15366 VSS.n8248 VSS.n8245 4.608
R15367 VSS.n8245 VSS.n8242 4.608
R15368 VSS.n8242 VSS.n8239 4.608
R15369 VSS.n8239 VSS.n8236 4.608
R15370 VSS.n8236 VSS.n8233 4.608
R15371 VSS.n8233 VSS.n8230 4.608
R15372 VSS.n8230 VSS.n8227 4.608
R15373 VSS.n8227 VSS.n8224 4.608
R15374 VSS.n8224 VSS.n8221 4.608
R15375 VSS.n8221 VSS.n8218 4.608
R15376 VSS.n8218 VSS.n8215 4.608
R15377 VSS.n8004 VSS.n8003 4.608
R15378 VSS.n8003 VSS.n8000 4.608
R15379 VSS.n8000 VSS.n7997 4.608
R15380 VSS.n7997 VSS.n7994 4.608
R15381 VSS.n7994 VSS.n7991 4.608
R15382 VSS.n7991 VSS.n7988 4.608
R15383 VSS.n7988 VSS.n7985 4.608
R15384 VSS.n7985 VSS.n7982 4.608
R15385 VSS.n7982 VSS.n7979 4.608
R15386 VSS.n7979 VSS.n7976 4.608
R15387 VSS.n7976 VSS.n7973 4.608
R15388 VSS.n7973 VSS.n7970 4.608
R15389 VSS.n7761 VSS.n7760 4.608
R15390 VSS.n7760 VSS.n7757 4.608
R15391 VSS.n7757 VSS.n7754 4.608
R15392 VSS.n7754 VSS.n7751 4.608
R15393 VSS.n7751 VSS.n7748 4.608
R15394 VSS.n7748 VSS.n7745 4.608
R15395 VSS.n7745 VSS.n7742 4.608
R15396 VSS.n7742 VSS.n7739 4.608
R15397 VSS.n7739 VSS.n7736 4.608
R15398 VSS.n7736 VSS.n7733 4.608
R15399 VSS.n7733 VSS.n7730 4.608
R15400 VSS.n7730 VSS.n7727 4.608
R15401 VSS.n7516 VSS.n7515 4.608
R15402 VSS.n7515 VSS.n7512 4.608
R15403 VSS.n7512 VSS.n7509 4.608
R15404 VSS.n7509 VSS.n7506 4.608
R15405 VSS.n7506 VSS.n7503 4.608
R15406 VSS.n7503 VSS.n7500 4.608
R15407 VSS.n7500 VSS.n7497 4.608
R15408 VSS.n7497 VSS.n7494 4.608
R15409 VSS.n7494 VSS.n7491 4.608
R15410 VSS.n7491 VSS.n7488 4.608
R15411 VSS.n7488 VSS.n7485 4.608
R15412 VSS.n7485 VSS.n7482 4.608
R15413 VSS.n1273 VSS.n1272 4.608
R15414 VSS.n1274 VSS.n1273 4.608
R15415 VSS.n1274 VSS.n646 4.608
R15416 VSS.n1280 VSS.n646 4.608
R15417 VSS.n1281 VSS.n1280 4.608
R15418 VSS.n1282 VSS.n1281 4.608
R15419 VSS.n1282 VSS.n642 4.608
R15420 VSS.n1288 VSS.n642 4.608
R15421 VSS.n1289 VSS.n1288 4.608
R15422 VSS.n1290 VSS.n1289 4.608
R15423 VSS.n1290 VSS.n638 4.608
R15424 VSS.n1296 VSS.n638 4.608
R15425 VSS.n914 VSS.n913 4.608
R15426 VSS.n913 VSS.n912 4.608
R15427 VSS.n912 VSS.n886 4.608
R15428 VSS.n906 VSS.n886 4.608
R15429 VSS.n906 VSS.n905 4.608
R15430 VSS.n905 VSS.n904 4.608
R15431 VSS.n904 VSS.n890 4.608
R15432 VSS.n898 VSS.n890 4.608
R15433 VSS.n898 VSS.n897 4.608
R15434 VSS.n897 VSS.n896 4.608
R15435 VSS.n896 VSS.n623 4.608
R15436 VSS.n1323 VSS.n623 4.608
R15437 VSS.n5700 VSS.n591 4.608
R15438 VSS.n5694 VSS.n591 4.608
R15439 VSS.n5694 VSS.n5693 4.608
R15440 VSS.n5693 VSS.n5692 4.608
R15441 VSS.n5692 VSS.n597 4.608
R15442 VSS.n5686 VSS.n597 4.608
R15443 VSS.n5686 VSS.n5685 4.608
R15444 VSS.n5685 VSS.n5684 4.608
R15445 VSS.n5684 VSS.n601 4.608
R15446 VSS.n5678 VSS.n601 4.608
R15447 VSS.n5678 VSS.n5677 4.608
R15448 VSS.n5677 VSS.n5676 4.608
R15449 VSS.n5619 VSS.n5618 4.608
R15450 VSS.n5619 VSS.n1376 4.608
R15451 VSS.n5625 VSS.n1376 4.608
R15452 VSS.n5626 VSS.n5625 4.608
R15453 VSS.n5627 VSS.n5626 4.608
R15454 VSS.n5627 VSS.n1372 4.608
R15455 VSS.n5633 VSS.n1372 4.608
R15456 VSS.n5634 VSS.n5633 4.608
R15457 VSS.n5636 VSS.n5634 4.608
R15458 VSS.n5636 VSS.n5635 4.608
R15459 VSS.n5635 VSS.n1368 4.608
R15460 VSS.n5643 VSS.n1368 4.608
R15461 VSS.n5492 VSS.n1448 4.608
R15462 VSS.n5486 VSS.n1448 4.608
R15463 VSS.n5486 VSS.n5485 4.608
R15464 VSS.n5485 VSS.n5484 4.608
R15465 VSS.n5484 VSS.n1452 4.608
R15466 VSS.n5478 VSS.n1452 4.608
R15467 VSS.n5478 VSS.n5477 4.608
R15468 VSS.n5477 VSS.n5476 4.608
R15469 VSS.n5476 VSS.n1456 4.608
R15470 VSS.n5470 VSS.n1456 4.608
R15471 VSS.n5470 VSS.n5469 4.608
R15472 VSS.n5469 VSS.n5468 4.608
R15473 VSS.n5411 VSS.n5410 4.608
R15474 VSS.n5411 VSS.n1517 4.608
R15475 VSS.n5417 VSS.n1517 4.608
R15476 VSS.n5418 VSS.n5417 4.608
R15477 VSS.n5419 VSS.n5418 4.608
R15478 VSS.n5419 VSS.n1513 4.608
R15479 VSS.n5425 VSS.n1513 4.608
R15480 VSS.n5426 VSS.n5425 4.608
R15481 VSS.n5428 VSS.n5426 4.608
R15482 VSS.n5428 VSS.n5427 4.608
R15483 VSS.n5427 VSS.n1509 4.608
R15484 VSS.n5435 VSS.n1509 4.608
R15485 VSS.n4759 VSS.n4727 4.608
R15486 VSS.n4753 VSS.n4727 4.608
R15487 VSS.n4753 VSS.n4752 4.608
R15488 VSS.n4752 VSS.n4751 4.608
R15489 VSS.n4751 VSS.n4731 4.608
R15490 VSS.n4745 VSS.n4731 4.608
R15491 VSS.n4745 VSS.n4744 4.608
R15492 VSS.n4744 VSS.n4743 4.608
R15493 VSS.n4743 VSS.n4735 4.608
R15494 VSS.n4737 VSS.n4735 4.608
R15495 VSS.n4737 VSS.n3124 4.608
R15496 VSS.n5079 VSS.n3124 4.608
R15497 VSS.n5023 VSS.n3151 4.608
R15498 VSS.n5029 VSS.n3151 4.608
R15499 VSS.n5030 VSS.n5029 4.608
R15500 VSS.n5031 VSS.n5030 4.608
R15501 VSS.n5031 VSS.n3147 4.608
R15502 VSS.n5037 VSS.n3147 4.608
R15503 VSS.n5038 VSS.n5037 4.608
R15504 VSS.n5039 VSS.n5038 4.608
R15505 VSS.n5039 VSS.n3143 4.608
R15506 VSS.n5045 VSS.n3143 4.608
R15507 VSS.n5046 VSS.n5045 4.608
R15508 VSS.n5047 VSS.n5046 4.608
R15509 VSS.n3232 VSS.n3220 4.608
R15510 VSS.n4524 VSS.n3232 4.608
R15511 VSS.n4524 VSS.n4523 4.608
R15512 VSS.n4523 VSS.n4522 4.608
R15513 VSS.n4522 VSS.n3233 4.608
R15514 VSS.n4516 VSS.n3233 4.608
R15515 VSS.n4516 VSS.n4515 4.608
R15516 VSS.n4515 VSS.n4514 4.608
R15517 VSS.n4514 VSS.n3237 4.608
R15518 VSS.n4508 VSS.n3237 4.608
R15519 VSS.n4508 VSS.n4507 4.608
R15520 VSS.n4507 VSS.n4506 4.608
R15521 VSS.n4169 VSS.n4137 4.608
R15522 VSS.n4163 VSS.n4137 4.608
R15523 VSS.n4163 VSS.n4162 4.608
R15524 VSS.n4162 VSS.n4161 4.608
R15525 VSS.n4161 VSS.n4141 4.608
R15526 VSS.n4155 VSS.n4141 4.608
R15527 VSS.n4155 VSS.n4154 4.608
R15528 VSS.n4154 VSS.n4153 4.608
R15529 VSS.n4153 VSS.n4145 4.608
R15530 VSS.n4147 VSS.n4145 4.608
R15531 VSS.n4147 VSS.n3294 4.608
R15532 VSS.n4475 VSS.n3294 4.608
R15533 VSS.n4424 VSS.n4423 4.608
R15534 VSS.n4425 VSS.n4424 4.608
R15535 VSS.n4425 VSS.n3316 4.608
R15536 VSS.n4431 VSS.n3316 4.608
R15537 VSS.n4432 VSS.n4431 4.608
R15538 VSS.n4433 VSS.n4432 4.608
R15539 VSS.n4433 VSS.n3312 4.608
R15540 VSS.n4439 VSS.n3312 4.608
R15541 VSS.n4440 VSS.n4439 4.608
R15542 VSS.n4441 VSS.n4440 4.608
R15543 VSS.n4441 VSS.n3308 4.608
R15544 VSS.n4447 VSS.n3308 4.608
R15545 VSS.n3950 VSS.n3392 4.608
R15546 VSS.n3396 VSS.n3392 4.608
R15547 VSS.n3943 VSS.n3396 4.608
R15548 VSS.n3943 VSS.n3942 4.608
R15549 VSS.n3942 VSS.n3941 4.608
R15550 VSS.n3941 VSS.n3397 4.608
R15551 VSS.n3935 VSS.n3397 4.608
R15552 VSS.n3935 VSS.n3934 4.608
R15553 VSS.n3934 VSS.n3933 4.608
R15554 VSS.n3933 VSS.n3401 4.608
R15555 VSS.n3927 VSS.n3401 4.608
R15556 VSS.n3927 VSS.n3926 4.608
R15557 VSS.n3557 VSS.n3525 4.608
R15558 VSS.n3551 VSS.n3525 4.608
R15559 VSS.n3551 VSS.n3550 4.608
R15560 VSS.n3550 VSS.n3549 4.608
R15561 VSS.n3549 VSS.n3529 4.608
R15562 VSS.n3543 VSS.n3529 4.608
R15563 VSS.n3543 VSS.n3542 4.608
R15564 VSS.n3542 VSS.n3541 4.608
R15565 VSS.n3541 VSS.n3533 4.608
R15566 VSS.n3535 VSS.n3533 4.608
R15567 VSS.n3535 VSS.n3420 4.608
R15568 VSS.n3864 VSS.n3420 4.608
R15569 VSS.n10564 VSS.n10563 4.589
R15570 VSS.n7082 VSS.n7081 4.524
R15571 VSS.n10566 VSS.n10565 4.5
R15572 VSS.n7045 VSS.n518 4.5
R15573 VSS.n7047 VSS.n7046 4.5
R15574 VSS.n496 VSS.n495 4.5
R15575 VSS.n495 VSS.n494 4.5
R15576 VSS VSS.n497 4.353
R15577 VSS.n16341 VSS.n16334 4.3
R15578 VSS.n16086 VSS.n16079 4.3
R15579 VSS.n15841 VSS.n15834 4.3
R15580 VSS.n15598 VSS.n15591 4.3
R15581 VSS.n15353 VSS.n15346 4.3
R15582 VSS.n15110 VSS.n15103 4.3
R15583 VSS.n14865 VSS.n14858 4.3
R15584 VSS.n12390 VSS.n12383 4.3
R15585 VSS.n12135 VSS.n12128 4.3
R15586 VSS.n11890 VSS.n11883 4.3
R15587 VSS.n11647 VSS.n11640 4.3
R15588 VSS.n11402 VSS.n11395 4.3
R15589 VSS.n11159 VSS.n11152 4.3
R15590 VSS.n10914 VSS.n10907 4.3
R15591 VSS.n8958 VSS.n8951 4.3
R15592 VSS.n8703 VSS.n8696 4.3
R15593 VSS.n8458 VSS.n8451 4.3
R15594 VSS.n8215 VSS.n8208 4.3
R15595 VSS.n7970 VSS.n7963 4.3
R15596 VSS.n7727 VSS.n7720 4.3
R15597 VSS.n7482 VSS.n7475 4.3
R15598 VSS.n1297 VSS.n1296 4.3
R15599 VSS.n1323 VSS.n1322 4.3
R15600 VSS.n5676 VSS.n605 4.3
R15601 VSS.n5644 VSS.n5643 4.3
R15602 VSS.n5468 VSS.n1460 4.3
R15603 VSS.n5436 VSS.n5435 4.3
R15604 VSS.n5080 VSS.n5079 4.3
R15605 VSS.n5047 VSS.n3138 4.3
R15606 VSS.n4506 VSS.n3241 4.3
R15607 VSS.n4475 VSS.n4474 4.3
R15608 VSS.n4448 VSS.n4447 4.3
R15609 VSS.n3926 VSS.n3925 4.3
R15610 VSS.n3865 VSS.n3864 4.3
R15611 VSS.n493 VSS.n492 4.235
R15612 VSS.n383 VSS.n370 4.141
R15613 VSS.n391 VSS.n368 4.141
R15614 VSS.n421 VSS.n350 4.141
R15615 VSS.n430 VSS.n347 4.141
R15616 VSS.n18175 VSS.n18162 4.141
R15617 VSS.n18183 VSS.n18160 4.141
R15618 VSS.n18215 VSS.n18142 4.141
R15619 VSS.n18220 VSS.n18140 4.141
R15620 VSS.n404 VSS.n362 4.137
R15621 VSS.n412 VSS.n357 4.137
R15622 VSS.n18196 VSS.n18154 4.137
R15623 VSS.n18204 VSS.n18149 4.137
R15624 VSS.n6939 VSS.n6938 4.116
R15625 VSS.n14478 VSS.n14477 4.088
R15626 VSS.n14298 VSS.n14297 4.088
R15627 VSS.n14491 VSS.n14490 4.088
R15628 VSS.n14503 VSS.n14502 4.088
R15629 VSS.n14515 VSS.n14514 4.088
R15630 VSS.n14527 VSS.n14526 4.088
R15631 VSS.n14539 VSS.n14538 4.088
R15632 VSS.n14551 VSS.n14550 4.088
R15633 VSS.n14076 VSS.n14075 4.088
R15634 VSS.n13895 VSS.n13894 4.088
R15635 VSS.n13715 VSS.n13714 4.088
R15636 VSS.n13535 VSS.n13534 4.088
R15637 VSS.n13355 VSS.n13354 4.088
R15638 VSS.n13175 VSS.n13174 4.088
R15639 VSS.n12995 VSS.n12994 4.088
R15640 VSS.n12815 VSS.n12814 4.088
R15641 VSS.n9219 VSS.n9218 4.088
R15642 VSS.n9387 VSS.n9386 4.088
R15643 VSS.n9555 VSS.n9554 4.088
R15644 VSS.n9723 VSS.n9722 4.088
R15645 VSS.n9891 VSS.n9890 4.088
R15646 VSS.n10059 VSS.n10058 4.088
R15647 VSS.n10227 VSS.n10226 4.088
R15648 VSS.n10394 VSS.n10393 4.088
R15649 VSS.n2462 VSS.n2461 4.088
R15650 VSS.n2552 VSS.n2551 4.088
R15651 VSS.n2642 VSS.n2641 4.088
R15652 VSS.n2732 VSS.n2731 4.088
R15653 VSS.n2822 VSS.n2821 4.088
R15654 VSS.n2912 VSS.n2911 4.088
R15655 VSS.n3002 VSS.n3001 4.088
R15656 VSS.n3092 VSS.n3091 4.088
R15657 VSS.n6240 VSS.n6239 4.088
R15658 VSS.n6304 VSS.n6303 4.088
R15659 VSS.n6368 VSS.n6367 4.088
R15660 VSS.n6383 VSS.n6382 4.088
R15661 VSS.n6936 VSS.n6935 4.088
R15662 VSS.n6846 VSS.n6845 4.088
R15663 VSS.n6756 VSS.n6755 4.088
R15664 VSS.n378 VSS.n375 4.019
R15665 VSS.n18170 VSS.n18167 4.019
R15666 VSS.n14643 VSS.n14642 4.008
R15667 VSS.n10692 VSS.n10691 4.008
R15668 VSS.n7260 VSS.n7259 4.008
R15669 VSS.n5134 VSS.n1654 4.008
R15670 VSS.n3451 VSS.n3446 4.008
R15671 VSS.n17532 VSS.n17531 3.732
R15672 VSS.n17364 VSS.n17363 3.732
R15673 VSS.n17196 VSS.n17195 3.732
R15674 VSS.n17028 VSS.n17027 3.732
R15675 VSS.n16860 VSS.n16859 3.732
R15676 VSS.n16692 VSS.n16691 3.732
R15677 VSS.n10497 VSS.n10496 3.732
R15678 VSS.n6248 VSS.n6077 3.732
R15679 VSS.n6312 VSS.n5961 3.732
R15680 VSS.n6376 VSS.n5845 3.732
R15681 VSS.n6941 VSS.n5789 3.732
R15682 VSS.n16609 VSS.n16608 3.582
R15683 VSS.n16621 VSS.n16620 3.582
R15684 VSS.n16636 VSS.n16635 3.582
R15685 VSS.n16645 VSS.n16644 3.582
R15686 VSS.n16657 VSS.n16656 3.582
R15687 VSS.n16669 VSS.n16668 3.582
R15688 VSS.n16681 VSS.n16680 3.582
R15689 VSS.n16740 VSS.n16739 3.582
R15690 VSS.n16777 VSS.n16776 3.582
R15691 VSS.n16789 VSS.n16788 3.582
R15692 VSS.n16804 VSS.n16803 3.582
R15693 VSS.n16813 VSS.n16812 3.582
R15694 VSS.n16825 VSS.n16824 3.582
R15695 VSS.n16837 VSS.n16836 3.582
R15696 VSS.n16849 VSS.n16848 3.582
R15697 VSS.n16908 VSS.n16907 3.582
R15698 VSS.n16945 VSS.n16944 3.582
R15699 VSS.n16957 VSS.n16956 3.582
R15700 VSS.n16972 VSS.n16971 3.582
R15701 VSS.n16981 VSS.n16980 3.582
R15702 VSS.n16993 VSS.n16992 3.582
R15703 VSS.n17005 VSS.n17004 3.582
R15704 VSS.n17017 VSS.n17016 3.582
R15705 VSS.n17076 VSS.n17075 3.582
R15706 VSS.n17113 VSS.n17112 3.582
R15707 VSS.n17125 VSS.n17124 3.582
R15708 VSS.n17140 VSS.n17139 3.582
R15709 VSS.n17149 VSS.n17148 3.582
R15710 VSS.n17161 VSS.n17160 3.582
R15711 VSS.n17173 VSS.n17172 3.582
R15712 VSS.n17185 VSS.n17184 3.582
R15713 VSS.n17244 VSS.n17243 3.582
R15714 VSS.n17281 VSS.n17280 3.582
R15715 VSS.n17293 VSS.n17292 3.582
R15716 VSS.n17308 VSS.n17307 3.582
R15717 VSS.n17317 VSS.n17316 3.582
R15718 VSS.n17329 VSS.n17328 3.582
R15719 VSS.n17341 VSS.n17340 3.582
R15720 VSS.n17353 VSS.n17352 3.582
R15721 VSS.n17412 VSS.n17411 3.582
R15722 VSS.n17449 VSS.n17448 3.582
R15723 VSS.n17461 VSS.n17460 3.582
R15724 VSS.n17476 VSS.n17475 3.582
R15725 VSS.n17485 VSS.n17484 3.582
R15726 VSS.n17497 VSS.n17496 3.582
R15727 VSS.n17509 VSS.n17508 3.582
R15728 VSS.n17521 VSS.n17520 3.582
R15729 VSS.n17580 VSS.n17579 3.582
R15730 VSS.n14223 VSS.n14222 3.582
R15731 VSS.n14211 VSS.n14210 3.582
R15732 VSS.n14199 VSS.n14198 3.582
R15733 VSS.n14187 VSS.n14186 3.582
R15734 VSS.n14175 VSS.n14174 3.582
R15735 VSS.n14163 VSS.n14162 3.582
R15736 VSS.n14151 VSS.n14150 3.582
R15737 VSS.n14139 VSS.n14138 3.582
R15738 VSS.n14403 VSS.n14402 3.582
R15739 VSS.n14391 VSS.n14390 3.582
R15740 VSS.n14379 VSS.n14378 3.582
R15741 VSS.n14367 VSS.n14366 3.582
R15742 VSS.n14355 VSS.n14354 3.582
R15743 VSS.n14343 VSS.n14342 3.582
R15744 VSS.n14331 VSS.n14330 3.582
R15745 VSS.n14319 VSS.n14318 3.582
R15746 VSS.n12740 VSS.n12739 3.582
R15747 VSS.n12728 VSS.n12727 3.582
R15748 VSS.n12716 VSS.n12715 3.582
R15749 VSS.n12704 VSS.n12703 3.582
R15750 VSS.n12692 VSS.n12691 3.582
R15751 VSS.n12680 VSS.n12679 3.582
R15752 VSS.n12668 VSS.n12667 3.582
R15753 VSS.n12656 VSS.n12655 3.582
R15754 VSS.n12920 VSS.n12919 3.582
R15755 VSS.n12908 VSS.n12907 3.582
R15756 VSS.n12896 VSS.n12895 3.582
R15757 VSS.n12884 VSS.n12883 3.582
R15758 VSS.n12872 VSS.n12871 3.582
R15759 VSS.n12860 VSS.n12859 3.582
R15760 VSS.n12848 VSS.n12847 3.582
R15761 VSS.n12836 VSS.n12835 3.582
R15762 VSS.n13100 VSS.n13099 3.582
R15763 VSS.n13088 VSS.n13087 3.582
R15764 VSS.n13076 VSS.n13075 3.582
R15765 VSS.n13064 VSS.n13063 3.582
R15766 VSS.n13052 VSS.n13051 3.582
R15767 VSS.n13040 VSS.n13039 3.582
R15768 VSS.n13028 VSS.n13027 3.582
R15769 VSS.n13016 VSS.n13015 3.582
R15770 VSS.n13280 VSS.n13279 3.582
R15771 VSS.n13268 VSS.n13267 3.582
R15772 VSS.n13256 VSS.n13255 3.582
R15773 VSS.n13244 VSS.n13243 3.582
R15774 VSS.n13232 VSS.n13231 3.582
R15775 VSS.n13220 VSS.n13219 3.582
R15776 VSS.n13208 VSS.n13207 3.582
R15777 VSS.n13196 VSS.n13195 3.582
R15778 VSS.n13460 VSS.n13459 3.582
R15779 VSS.n13448 VSS.n13447 3.582
R15780 VSS.n13436 VSS.n13435 3.582
R15781 VSS.n13424 VSS.n13423 3.582
R15782 VSS.n13412 VSS.n13411 3.582
R15783 VSS.n13400 VSS.n13399 3.582
R15784 VSS.n13388 VSS.n13387 3.582
R15785 VSS.n13376 VSS.n13375 3.582
R15786 VSS.n13640 VSS.n13639 3.582
R15787 VSS.n13628 VSS.n13627 3.582
R15788 VSS.n13616 VSS.n13615 3.582
R15789 VSS.n13604 VSS.n13603 3.582
R15790 VSS.n13592 VSS.n13591 3.582
R15791 VSS.n13580 VSS.n13579 3.582
R15792 VSS.n13568 VSS.n13567 3.582
R15793 VSS.n13556 VSS.n13555 3.582
R15794 VSS.n13820 VSS.n13819 3.582
R15795 VSS.n13808 VSS.n13807 3.582
R15796 VSS.n13796 VSS.n13795 3.582
R15797 VSS.n13784 VSS.n13783 3.582
R15798 VSS.n13772 VSS.n13771 3.582
R15799 VSS.n13760 VSS.n13759 3.582
R15800 VSS.n13748 VSS.n13747 3.582
R15801 VSS.n13736 VSS.n13735 3.582
R15802 VSS.n14000 VSS.n13999 3.582
R15803 VSS.n13988 VSS.n13987 3.582
R15804 VSS.n13976 VSS.n13975 3.582
R15805 VSS.n13964 VSS.n13963 3.582
R15806 VSS.n13952 VSS.n13951 3.582
R15807 VSS.n13940 VSS.n13939 3.582
R15808 VSS.n13928 VSS.n13927 3.582
R15809 VSS.n13916 VSS.n13915 3.582
R15810 VSS.n10247 VSS.n10246 3.582
R15811 VSS.n10259 VSS.n10258 3.582
R15812 VSS.n10274 VSS.n10273 3.582
R15813 VSS.n10283 VSS.n10282 3.582
R15814 VSS.n10295 VSS.n10294 3.582
R15815 VSS.n10307 VSS.n10306 3.582
R15816 VSS.n10319 VSS.n10318 3.582
R15817 VSS.n10376 VSS.n10375 3.582
R15818 VSS.n10079 VSS.n10078 3.582
R15819 VSS.n10091 VSS.n10090 3.582
R15820 VSS.n10106 VSS.n10105 3.582
R15821 VSS.n10115 VSS.n10114 3.582
R15822 VSS.n10127 VSS.n10126 3.582
R15823 VSS.n10139 VSS.n10138 3.582
R15824 VSS.n10151 VSS.n10150 3.582
R15825 VSS.n10208 VSS.n10207 3.582
R15826 VSS.n9911 VSS.n9910 3.582
R15827 VSS.n9923 VSS.n9922 3.582
R15828 VSS.n9938 VSS.n9937 3.582
R15829 VSS.n9947 VSS.n9946 3.582
R15830 VSS.n9959 VSS.n9958 3.582
R15831 VSS.n9971 VSS.n9970 3.582
R15832 VSS.n9983 VSS.n9982 3.582
R15833 VSS.n10040 VSS.n10039 3.582
R15834 VSS.n9743 VSS.n9742 3.582
R15835 VSS.n9755 VSS.n9754 3.582
R15836 VSS.n9770 VSS.n9769 3.582
R15837 VSS.n9779 VSS.n9778 3.582
R15838 VSS.n9791 VSS.n9790 3.582
R15839 VSS.n9803 VSS.n9802 3.582
R15840 VSS.n9815 VSS.n9814 3.582
R15841 VSS.n9872 VSS.n9871 3.582
R15842 VSS.n9575 VSS.n9574 3.582
R15843 VSS.n9587 VSS.n9586 3.582
R15844 VSS.n9602 VSS.n9601 3.582
R15845 VSS.n9611 VSS.n9610 3.582
R15846 VSS.n9623 VSS.n9622 3.582
R15847 VSS.n9635 VSS.n9634 3.582
R15848 VSS.n9647 VSS.n9646 3.582
R15849 VSS.n9704 VSS.n9703 3.582
R15850 VSS.n9407 VSS.n9406 3.582
R15851 VSS.n9419 VSS.n9418 3.582
R15852 VSS.n9434 VSS.n9433 3.582
R15853 VSS.n9443 VSS.n9442 3.582
R15854 VSS.n9455 VSS.n9454 3.582
R15855 VSS.n9467 VSS.n9466 3.582
R15856 VSS.n9479 VSS.n9478 3.582
R15857 VSS.n9536 VSS.n9535 3.582
R15858 VSS.n9239 VSS.n9238 3.582
R15859 VSS.n9251 VSS.n9250 3.582
R15860 VSS.n9266 VSS.n9265 3.582
R15861 VSS.n9275 VSS.n9274 3.582
R15862 VSS.n9287 VSS.n9286 3.582
R15863 VSS.n9299 VSS.n9298 3.582
R15864 VSS.n9311 VSS.n9310 3.582
R15865 VSS.n9368 VSS.n9367 3.582
R15866 VSS.n10426 VSS.n10425 3.582
R15867 VSS.n10450 VSS.n10449 3.582
R15868 VSS.n10474 VSS.n10473 3.582
R15869 VSS.n10544 VSS.n10543 3.582
R15870 VSS.n10486 VSS.n10485 3.582
R15871 VSS.n10462 VSS.n10461 3.582
R15872 VSS.n10441 VSS.n10440 3.582
R15873 VSS.n10414 VSS.n10413 3.582
R15874 VSS.n1689 VSS.n1683 3.582
R15875 VSS.n3055 VSS.n1690 3.582
R15876 VSS.n3061 VSS.n1691 3.582
R15877 VSS.n3067 VSS.n1687 3.582
R15878 VSS.n3073 VSS.n1692 3.582
R15879 VSS.n3082 VSS.n1686 3.582
R15880 VSS.n3087 VSS.n1693 3.582
R15881 VSS.n1779 VSS.n1773 3.582
R15882 VSS.n2965 VSS.n1780 3.582
R15883 VSS.n2971 VSS.n1781 3.582
R15884 VSS.n2977 VSS.n1777 3.582
R15885 VSS.n2983 VSS.n1782 3.582
R15886 VSS.n2992 VSS.n1776 3.582
R15887 VSS.n2997 VSS.n1783 3.582
R15888 VSS.n1869 VSS.n1863 3.582
R15889 VSS.n2875 VSS.n1870 3.582
R15890 VSS.n2881 VSS.n1871 3.582
R15891 VSS.n2887 VSS.n1867 3.582
R15892 VSS.n2893 VSS.n1872 3.582
R15893 VSS.n2902 VSS.n1866 3.582
R15894 VSS.n2907 VSS.n1873 3.582
R15895 VSS.n1959 VSS.n1953 3.582
R15896 VSS.n2785 VSS.n1960 3.582
R15897 VSS.n2791 VSS.n1961 3.582
R15898 VSS.n2797 VSS.n1957 3.582
R15899 VSS.n2803 VSS.n1962 3.582
R15900 VSS.n2812 VSS.n1956 3.582
R15901 VSS.n2817 VSS.n1963 3.582
R15902 VSS.n2049 VSS.n2043 3.582
R15903 VSS.n2695 VSS.n2050 3.582
R15904 VSS.n2701 VSS.n2051 3.582
R15905 VSS.n2707 VSS.n2047 3.582
R15906 VSS.n2713 VSS.n2052 3.582
R15907 VSS.n2722 VSS.n2046 3.582
R15908 VSS.n2727 VSS.n2053 3.582
R15909 VSS.n2139 VSS.n2133 3.582
R15910 VSS.n2605 VSS.n2140 3.582
R15911 VSS.n2611 VSS.n2141 3.582
R15912 VSS.n2617 VSS.n2137 3.582
R15913 VSS.n2623 VSS.n2142 3.582
R15914 VSS.n2632 VSS.n2136 3.582
R15915 VSS.n2637 VSS.n2143 3.582
R15916 VSS.n2229 VSS.n2223 3.582
R15917 VSS.n2515 VSS.n2230 3.582
R15918 VSS.n2521 VSS.n2231 3.582
R15919 VSS.n2527 VSS.n2227 3.582
R15920 VSS.n2533 VSS.n2232 3.582
R15921 VSS.n2542 VSS.n2226 3.582
R15922 VSS.n2547 VSS.n2233 3.582
R15923 VSS.n2319 VSS.n2313 3.582
R15924 VSS.n2425 VSS.n2320 3.582
R15925 VSS.n2431 VSS.n2321 3.582
R15926 VSS.n2437 VSS.n2317 3.582
R15927 VSS.n2443 VSS.n2322 3.582
R15928 VSS.n2452 VSS.n2316 3.582
R15929 VSS.n2457 VSS.n2323 3.582
R15930 VSS.n2414 VSS.n2318 3.582
R15931 VSS.n2504 VSS.n2228 3.582
R15932 VSS.n2594 VSS.n2138 3.582
R15933 VSS.n2684 VSS.n2048 3.582
R15934 VSS.n2774 VSS.n1958 3.582
R15935 VSS.n2864 VSS.n1868 3.582
R15936 VSS.n2954 VSS.n1778 3.582
R15937 VSS.n3044 VSS.n1688 3.582
R15938 VSS.n6613 VSS.n6607 3.582
R15939 VSS.n6712 VSS.n6614 3.582
R15940 VSS.n6718 VSS.n6612 3.582
R15941 VSS.n6724 VSS.n6615 3.582
R15942 VSS.n6730 VSS.n6611 3.582
R15943 VSS.n6736 VSS.n6616 3.582
R15944 VSS.n6745 VSS.n6610 3.582
R15945 VSS.n6750 VSS.n6617 3.582
R15946 VSS.n6523 VSS.n6517 3.582
R15947 VSS.n6802 VSS.n6524 3.582
R15948 VSS.n6808 VSS.n6522 3.582
R15949 VSS.n6814 VSS.n6525 3.582
R15950 VSS.n6820 VSS.n6521 3.582
R15951 VSS.n6826 VSS.n6526 3.582
R15952 VSS.n6835 VSS.n6520 3.582
R15953 VSS.n6840 VSS.n6527 3.582
R15954 VSS.n6433 VSS.n6427 3.582
R15955 VSS.n6892 VSS.n6434 3.582
R15956 VSS.n6898 VSS.n6432 3.582
R15957 VSS.n6904 VSS.n6435 3.582
R15958 VSS.n6910 VSS.n6431 3.582
R15959 VSS.n6916 VSS.n6436 3.582
R15960 VSS.n6925 VSS.n6430 3.582
R15961 VSS.n6930 VSS.n6437 3.582
R15962 VSS.n6174 VSS.n6099 3.582
R15963 VSS.n6158 VSS.n6106 3.582
R15964 VSS.n6142 VSS.n6100 3.582
R15965 VSS.n6126 VSS.n6105 3.582
R15966 VSS.n6134 VSS.n6104 3.582
R15967 VSS.n6150 VSS.n6101 3.582
R15968 VSS.n6166 VSS.n6103 3.582
R15969 VSS.n6182 VSS.n6102 3.582
R15970 VSS.n6058 VSS.n5983 3.582
R15971 VSS.n6042 VSS.n5990 3.582
R15972 VSS.n6026 VSS.n5984 3.582
R15973 VSS.n6010 VSS.n5989 3.582
R15974 VSS.n6018 VSS.n5988 3.582
R15975 VSS.n6034 VSS.n5985 3.582
R15976 VSS.n6050 VSS.n5987 3.582
R15977 VSS.n6066 VSS.n5986 3.582
R15978 VSS.n5942 VSS.n5867 3.582
R15979 VSS.n5926 VSS.n5874 3.582
R15980 VSS.n5910 VSS.n5868 3.582
R15981 VSS.n5894 VSS.n5873 3.582
R15982 VSS.n5902 VSS.n5872 3.582
R15983 VSS.n5918 VSS.n5869 3.582
R15984 VSS.n5934 VSS.n5871 3.582
R15985 VSS.n5950 VSS.n5870 3.582
R15986 VSS.n7006 VSS.n7005 3.582
R15987 VSS.n7018 VSS.n7017 3.582
R15988 VSS.n7030 VSS.n7029 3.582
R15989 VSS.n7042 VSS.n7041 3.582
R15990 VSS.n7036 VSS.n7035 3.582
R15991 VSS.n7024 VSS.n7023 3.582
R15992 VSS.n7012 VSS.n7011 3.582
R15993 VSS.n7000 VSS.n6999 3.582
R15994 VSS.t78 VSS.n17924 3.486
R15995 VSS.n17768 VSS.n17742 3.455
R15996 VSS.n17743 VSS.n17742 3.412
R15997 VSS.n377 VSS.n374 3.388
R15998 VSS.n384 VSS.n372 3.388
R15999 VSS.n429 VSS.n348 3.388
R16000 VSS.n435 VSS.n434 3.388
R16001 VSS.n18169 VSS.n18166 3.388
R16002 VSS.n18176 VSS.n18164 3.388
R16003 VSS.n18221 VSS.n18137 3.388
R16004 VSS.n18227 VSS.n18226 3.388
R16005 VSS VSS.n18026 3.308
R16006 VSS.n471 VSS 3.035
R16007 VSS.n7060 VSS 3.031
R16008 VSS.n17985 VSS 3.022
R16009 VSS.n380 VSS.n374 3.011
R16010 VSS.n380 VSS.n372 3.011
R16011 VSS.n348 VSS.n345 3.011
R16012 VSS.n434 VSS.n345 3.011
R16013 VSS.n18172 VSS.n18166 3.011
R16014 VSS.n18172 VSS.n18164 3.011
R16015 VSS.n18225 VSS.n18137 3.011
R16016 VSS.n18226 VSS.n18225 3.011
R16017 VSS.n16378 VSS.n16377 2.917
R16018 VSS.n16122 VSS.n16121 2.917
R16019 VSS.n15878 VSS.n15877 2.917
R16020 VSS.n15634 VSS.n15633 2.917
R16021 VSS.n15390 VSS.n15389 2.917
R16022 VSS.n15146 VSS.n15145 2.917
R16023 VSS.n14902 VSS.n14901 2.917
R16024 VSS.n12427 VSS.n12426 2.917
R16025 VSS.n12171 VSS.n12170 2.917
R16026 VSS.n11927 VSS.n11926 2.917
R16027 VSS.n11683 VSS.n11682 2.917
R16028 VSS.n11439 VSS.n11438 2.917
R16029 VSS.n11195 VSS.n11194 2.917
R16030 VSS.n10951 VSS.n10950 2.917
R16031 VSS.n8995 VSS.n8994 2.917
R16032 VSS.n8739 VSS.n8738 2.917
R16033 VSS.n8495 VSS.n8494 2.917
R16034 VSS.n8251 VSS.n8250 2.917
R16035 VSS.n8007 VSS.n8006 2.917
R16036 VSS.n7763 VSS.n7762 2.917
R16037 VSS.n7519 VSS.n7518 2.917
R16038 VSS.n4928 VSS.n4760 2.917
R16039 VSS.n5022 VSS.n5021 2.917
R16040 VSS.n4544 VSS.n4543 2.917
R16041 VSS.n4319 VSS.n4170 2.917
R16042 VSS.n4412 VSS.n3320 2.917
R16043 VSS.n3951 VSS.n3382 2.917
R16044 VSS.n3715 VSS.n3558 2.917
R16045 VSS.n1261 VSS.n650 2.917
R16046 VSS.n885 VSS.n712 2.917
R16047 VSS.n5701 VSS.n589 2.917
R16048 VSS.n5617 VSS.n1381 2.917
R16049 VSS.n5493 VSS.n1447 2.917
R16050 VSS.n5409 VSS.n1522 2.917
R16051 VSS.n482 VSS.t212 2.721
R16052 VSS.n16377 VSS.n16376 2.715
R16053 VSS.n16121 VSS.n16044 2.715
R16054 VSS.n15877 VSS.n15876 2.715
R16055 VSS.n15633 VSS.n15556 2.715
R16056 VSS.n15389 VSS.n15388 2.715
R16057 VSS.n15145 VSS.n15068 2.715
R16058 VSS.n14901 VSS.n14900 2.715
R16059 VSS.n12426 VSS.n12425 2.715
R16060 VSS.n12170 VSS.n12093 2.715
R16061 VSS.n11926 VSS.n11925 2.715
R16062 VSS.n11682 VSS.n11605 2.715
R16063 VSS.n11438 VSS.n11437 2.715
R16064 VSS.n11194 VSS.n11117 2.715
R16065 VSS.n10950 VSS.n10949 2.715
R16066 VSS.n8994 VSS.n8993 2.715
R16067 VSS.n8738 VSS.n8661 2.715
R16068 VSS.n8494 VSS.n8493 2.715
R16069 VSS.n8250 VSS.n8173 2.715
R16070 VSS.n8006 VSS.n8005 2.715
R16071 VSS.n7762 VSS.n7685 2.715
R16072 VSS.n7518 VSS.n7517 2.715
R16073 VSS.n1262 VSS.n650 2.715
R16074 VSS.n885 VSS.n884 2.715
R16075 VSS.n5702 VSS.n5701 2.715
R16076 VSS.n5617 VSS.n5616 2.715
R16077 VSS.n5493 VSS.n1446 2.715
R16078 VSS.n5409 VSS.n5408 2.715
R16079 VSS.n4760 VSS.n4726 2.715
R16080 VSS.n5022 VSS.n3156 2.715
R16081 VSS.n4543 VSS.n4542 2.715
R16082 VSS.n4170 VSS.n4136 2.715
R16083 VSS.n4413 VSS.n3320 2.715
R16084 VSS.n3952 VSS.n3951 2.715
R16085 VSS.n3558 VSS.n3524 2.715
R16086 VSS.n18021 VSS.n18020 2.554
R16087 VSS.n18230 VSS.n18229 2.529
R16088 VSS.n17948 VSS.n17923 2.488
R16089 VSS VSS.n18231 2.44
R16090 VSS.n439 VSS 2.37
R16091 VSS.n14077 VSS.n14076 2.287
R16092 VSS.n14097 VSS.n14084 2.26
R16093 VSS.n387 VSS.n370 2.258
R16094 VSS.n387 VSS.n368 2.258
R16095 VSS.n425 VSS.n350 2.258
R16096 VSS.n425 VSS.n347 2.258
R16097 VSS.n18179 VSS.n18162 2.258
R16098 VSS.n18179 VSS.n18160 2.258
R16099 VSS.n18216 VSS.n18215 2.258
R16100 VSS.n18216 VSS.n18140 2.258
R16101 VSS.n14082 VSS.n14081 2.245
R16102 VSS.n493 VSS.n472 2.241
R16103 VSS.n14098 VSS.n14083 2.239
R16104 VSS.n376 VSS.n375 2.228
R16105 VSS.n18168 VSS.n18167 2.228
R16106 VSS.n14649 VSS.n14648 1.95
R16107 VSS.n10698 VSS.n10697 1.95
R16108 VSS.n7266 VSS.n7265 1.95
R16109 VSS.n1653 VSS.n1586 1.95
R16110 VSS.n3448 VSS.n3447 1.95
R16111 VSS.n17807 VSS.n17806 1.95
R16112 VSS.n14079 VSS.n14078 1.901
R16113 VSS.n18327 VSS.n0 1.874
R16114 VSS.n260 VSS.n259 1.874
R16115 VSS.n14320 VSS.n14315 1.777
R16116 VSS.n14322 VSS.n14320 1.777
R16117 VSS.n14332 VSS.n14327 1.777
R16118 VSS.n14334 VSS.n14332 1.777
R16119 VSS.n14344 VSS.n14339 1.777
R16120 VSS.n14346 VSS.n14344 1.777
R16121 VSS.n14356 VSS.n14351 1.777
R16122 VSS.n14358 VSS.n14356 1.777
R16123 VSS.n14368 VSS.n14363 1.777
R16124 VSS.n14370 VSS.n14368 1.777
R16125 VSS.n14380 VSS.n14375 1.777
R16126 VSS.n14392 VSS.n14387 1.777
R16127 VSS.n14394 VSS.n14392 1.777
R16128 VSS.n14404 VSS.n14399 1.777
R16129 VSS.n14406 VSS.n14404 1.777
R16130 VSS.n14461 VSS.n14411 1.777
R16131 VSS.n14463 VSS.n14461 1.777
R16132 VSS.n14140 VSS.n14135 1.777
R16133 VSS.n14142 VSS.n14140 1.777
R16134 VSS.n14152 VSS.n14147 1.777
R16135 VSS.n14154 VSS.n14152 1.777
R16136 VSS.n14164 VSS.n14159 1.777
R16137 VSS.n14166 VSS.n14164 1.777
R16138 VSS.n14176 VSS.n14171 1.777
R16139 VSS.n14178 VSS.n14176 1.777
R16140 VSS.n14188 VSS.n14183 1.777
R16141 VSS.n14190 VSS.n14188 1.777
R16142 VSS.n14200 VSS.n14195 1.777
R16143 VSS.n14212 VSS.n14207 1.777
R16144 VSS.n14214 VSS.n14212 1.777
R16145 VSS.n14224 VSS.n14219 1.777
R16146 VSS.n14226 VSS.n14224 1.777
R16147 VSS.n14281 VSS.n14231 1.777
R16148 VSS.n14283 VSS.n14281 1.777
R16149 VSS.n17581 VSS.n17529 1.777
R16150 VSS.n17583 VSS.n17581 1.777
R16151 VSS.n17522 VSS.n17517 1.777
R16152 VSS.n17524 VSS.n17522 1.777
R16153 VSS.n17510 VSS.n17505 1.777
R16154 VSS.n17512 VSS.n17510 1.777
R16155 VSS.n17498 VSS.n17493 1.777
R16156 VSS.n17500 VSS.n17498 1.777
R16157 VSS.n17486 VSS.n17481 1.777
R16158 VSS.n17488 VSS.n17486 1.777
R16159 VSS.n17477 VSS.n17470 1.777
R16160 VSS.n17462 VSS.n17457 1.777
R16161 VSS.n17464 VSS.n17462 1.777
R16162 VSS.n17450 VSS.n17445 1.777
R16163 VSS.n17452 VSS.n17450 1.777
R16164 VSS.n17438 VSS.n17433 1.777
R16165 VSS.n17440 VSS.n17438 1.777
R16166 VSS.n17413 VSS.n17361 1.777
R16167 VSS.n17415 VSS.n17413 1.777
R16168 VSS.n17354 VSS.n17349 1.777
R16169 VSS.n17356 VSS.n17354 1.777
R16170 VSS.n17342 VSS.n17337 1.777
R16171 VSS.n17344 VSS.n17342 1.777
R16172 VSS.n17330 VSS.n17325 1.777
R16173 VSS.n17332 VSS.n17330 1.777
R16174 VSS.n17318 VSS.n17313 1.777
R16175 VSS.n17320 VSS.n17318 1.777
R16176 VSS.n17309 VSS.n17302 1.777
R16177 VSS.n17294 VSS.n17289 1.777
R16178 VSS.n17296 VSS.n17294 1.777
R16179 VSS.n17282 VSS.n17277 1.777
R16180 VSS.n17284 VSS.n17282 1.777
R16181 VSS.n17270 VSS.n17265 1.777
R16182 VSS.n17272 VSS.n17270 1.777
R16183 VSS.n17245 VSS.n17193 1.777
R16184 VSS.n17247 VSS.n17245 1.777
R16185 VSS.n17186 VSS.n17181 1.777
R16186 VSS.n17188 VSS.n17186 1.777
R16187 VSS.n17174 VSS.n17169 1.777
R16188 VSS.n17176 VSS.n17174 1.777
R16189 VSS.n17162 VSS.n17157 1.777
R16190 VSS.n17164 VSS.n17162 1.777
R16191 VSS.n17150 VSS.n17145 1.777
R16192 VSS.n17152 VSS.n17150 1.777
R16193 VSS.n17141 VSS.n17134 1.777
R16194 VSS.n17126 VSS.n17121 1.777
R16195 VSS.n17128 VSS.n17126 1.777
R16196 VSS.n17114 VSS.n17109 1.777
R16197 VSS.n17116 VSS.n17114 1.777
R16198 VSS.n17102 VSS.n17097 1.777
R16199 VSS.n17104 VSS.n17102 1.777
R16200 VSS.n17077 VSS.n17025 1.777
R16201 VSS.n17079 VSS.n17077 1.777
R16202 VSS.n17018 VSS.n17013 1.777
R16203 VSS.n17020 VSS.n17018 1.777
R16204 VSS.n17006 VSS.n17001 1.777
R16205 VSS.n17008 VSS.n17006 1.777
R16206 VSS.n16994 VSS.n16989 1.777
R16207 VSS.n16996 VSS.n16994 1.777
R16208 VSS.n16982 VSS.n16977 1.777
R16209 VSS.n16984 VSS.n16982 1.777
R16210 VSS.n16973 VSS.n16966 1.777
R16211 VSS.n16958 VSS.n16953 1.777
R16212 VSS.n16960 VSS.n16958 1.777
R16213 VSS.n16946 VSS.n16941 1.777
R16214 VSS.n16948 VSS.n16946 1.777
R16215 VSS.n16934 VSS.n16929 1.777
R16216 VSS.n16936 VSS.n16934 1.777
R16217 VSS.n16909 VSS.n16857 1.777
R16218 VSS.n16911 VSS.n16909 1.777
R16219 VSS.n16850 VSS.n16845 1.777
R16220 VSS.n16852 VSS.n16850 1.777
R16221 VSS.n16838 VSS.n16833 1.777
R16222 VSS.n16840 VSS.n16838 1.777
R16223 VSS.n16826 VSS.n16821 1.777
R16224 VSS.n16828 VSS.n16826 1.777
R16225 VSS.n16814 VSS.n16809 1.777
R16226 VSS.n16816 VSS.n16814 1.777
R16227 VSS.n16805 VSS.n16798 1.777
R16228 VSS.n16790 VSS.n16785 1.777
R16229 VSS.n16792 VSS.n16790 1.777
R16230 VSS.n16778 VSS.n16773 1.777
R16231 VSS.n16780 VSS.n16778 1.777
R16232 VSS.n16766 VSS.n16761 1.777
R16233 VSS.n16768 VSS.n16766 1.777
R16234 VSS.n16741 VSS.n16689 1.777
R16235 VSS.n16743 VSS.n16741 1.777
R16236 VSS.n16682 VSS.n16677 1.777
R16237 VSS.n16684 VSS.n16682 1.777
R16238 VSS.n16670 VSS.n16665 1.777
R16239 VSS.n16672 VSS.n16670 1.777
R16240 VSS.n16658 VSS.n16653 1.777
R16241 VSS.n16660 VSS.n16658 1.777
R16242 VSS.n16646 VSS.n16641 1.777
R16243 VSS.n16648 VSS.n16646 1.777
R16244 VSS.n16637 VSS.n16630 1.777
R16245 VSS.n16622 VSS.n16617 1.777
R16246 VSS.n16624 VSS.n16622 1.777
R16247 VSS.n16610 VSS.n16605 1.777
R16248 VSS.n16612 VSS.n16610 1.777
R16249 VSS.n16598 VSS.n16593 1.777
R16250 VSS.n16600 VSS.n16598 1.777
R16251 VSS.n13917 VSS.n13912 1.777
R16252 VSS.n13919 VSS.n13917 1.777
R16253 VSS.n13929 VSS.n13924 1.777
R16254 VSS.n13931 VSS.n13929 1.777
R16255 VSS.n13941 VSS.n13936 1.777
R16256 VSS.n13943 VSS.n13941 1.777
R16257 VSS.n13953 VSS.n13948 1.777
R16258 VSS.n13955 VSS.n13953 1.777
R16259 VSS.n13965 VSS.n13960 1.777
R16260 VSS.n13967 VSS.n13965 1.777
R16261 VSS.n13977 VSS.n13972 1.777
R16262 VSS.n13989 VSS.n13984 1.777
R16263 VSS.n13991 VSS.n13989 1.777
R16264 VSS.n14001 VSS.n13996 1.777
R16265 VSS.n14003 VSS.n14001 1.777
R16266 VSS.n14058 VSS.n14008 1.777
R16267 VSS.n14060 VSS.n14058 1.777
R16268 VSS.n13737 VSS.n13732 1.777
R16269 VSS.n13739 VSS.n13737 1.777
R16270 VSS.n13749 VSS.n13744 1.777
R16271 VSS.n13751 VSS.n13749 1.777
R16272 VSS.n13761 VSS.n13756 1.777
R16273 VSS.n13763 VSS.n13761 1.777
R16274 VSS.n13773 VSS.n13768 1.777
R16275 VSS.n13775 VSS.n13773 1.777
R16276 VSS.n13785 VSS.n13780 1.777
R16277 VSS.n13787 VSS.n13785 1.777
R16278 VSS.n13797 VSS.n13792 1.777
R16279 VSS.n13809 VSS.n13804 1.777
R16280 VSS.n13811 VSS.n13809 1.777
R16281 VSS.n13821 VSS.n13816 1.777
R16282 VSS.n13823 VSS.n13821 1.777
R16283 VSS.n13878 VSS.n13828 1.777
R16284 VSS.n13880 VSS.n13878 1.777
R16285 VSS.n13557 VSS.n13552 1.777
R16286 VSS.n13559 VSS.n13557 1.777
R16287 VSS.n13569 VSS.n13564 1.777
R16288 VSS.n13571 VSS.n13569 1.777
R16289 VSS.n13581 VSS.n13576 1.777
R16290 VSS.n13583 VSS.n13581 1.777
R16291 VSS.n13593 VSS.n13588 1.777
R16292 VSS.n13595 VSS.n13593 1.777
R16293 VSS.n13605 VSS.n13600 1.777
R16294 VSS.n13607 VSS.n13605 1.777
R16295 VSS.n13617 VSS.n13612 1.777
R16296 VSS.n13629 VSS.n13624 1.777
R16297 VSS.n13631 VSS.n13629 1.777
R16298 VSS.n13641 VSS.n13636 1.777
R16299 VSS.n13643 VSS.n13641 1.777
R16300 VSS.n13698 VSS.n13648 1.777
R16301 VSS.n13700 VSS.n13698 1.777
R16302 VSS.n13377 VSS.n13372 1.777
R16303 VSS.n13379 VSS.n13377 1.777
R16304 VSS.n13389 VSS.n13384 1.777
R16305 VSS.n13391 VSS.n13389 1.777
R16306 VSS.n13401 VSS.n13396 1.777
R16307 VSS.n13403 VSS.n13401 1.777
R16308 VSS.n13413 VSS.n13408 1.777
R16309 VSS.n13415 VSS.n13413 1.777
R16310 VSS.n13425 VSS.n13420 1.777
R16311 VSS.n13427 VSS.n13425 1.777
R16312 VSS.n13437 VSS.n13432 1.777
R16313 VSS.n13449 VSS.n13444 1.777
R16314 VSS.n13451 VSS.n13449 1.777
R16315 VSS.n13461 VSS.n13456 1.777
R16316 VSS.n13463 VSS.n13461 1.777
R16317 VSS.n13518 VSS.n13468 1.777
R16318 VSS.n13520 VSS.n13518 1.777
R16319 VSS.n13197 VSS.n13192 1.777
R16320 VSS.n13199 VSS.n13197 1.777
R16321 VSS.n13209 VSS.n13204 1.777
R16322 VSS.n13211 VSS.n13209 1.777
R16323 VSS.n13221 VSS.n13216 1.777
R16324 VSS.n13223 VSS.n13221 1.777
R16325 VSS.n13233 VSS.n13228 1.777
R16326 VSS.n13235 VSS.n13233 1.777
R16327 VSS.n13245 VSS.n13240 1.777
R16328 VSS.n13247 VSS.n13245 1.777
R16329 VSS.n13257 VSS.n13252 1.777
R16330 VSS.n13269 VSS.n13264 1.777
R16331 VSS.n13271 VSS.n13269 1.777
R16332 VSS.n13281 VSS.n13276 1.777
R16333 VSS.n13283 VSS.n13281 1.777
R16334 VSS.n13338 VSS.n13288 1.777
R16335 VSS.n13340 VSS.n13338 1.777
R16336 VSS.n13017 VSS.n13012 1.777
R16337 VSS.n13019 VSS.n13017 1.777
R16338 VSS.n13029 VSS.n13024 1.777
R16339 VSS.n13031 VSS.n13029 1.777
R16340 VSS.n13041 VSS.n13036 1.777
R16341 VSS.n13043 VSS.n13041 1.777
R16342 VSS.n13053 VSS.n13048 1.777
R16343 VSS.n13055 VSS.n13053 1.777
R16344 VSS.n13065 VSS.n13060 1.777
R16345 VSS.n13067 VSS.n13065 1.777
R16346 VSS.n13077 VSS.n13072 1.777
R16347 VSS.n13089 VSS.n13084 1.777
R16348 VSS.n13091 VSS.n13089 1.777
R16349 VSS.n13101 VSS.n13096 1.777
R16350 VSS.n13103 VSS.n13101 1.777
R16351 VSS.n13158 VSS.n13108 1.777
R16352 VSS.n13160 VSS.n13158 1.777
R16353 VSS.n12837 VSS.n12832 1.777
R16354 VSS.n12839 VSS.n12837 1.777
R16355 VSS.n12849 VSS.n12844 1.777
R16356 VSS.n12851 VSS.n12849 1.777
R16357 VSS.n12861 VSS.n12856 1.777
R16358 VSS.n12863 VSS.n12861 1.777
R16359 VSS.n12873 VSS.n12868 1.777
R16360 VSS.n12875 VSS.n12873 1.777
R16361 VSS.n12885 VSS.n12880 1.777
R16362 VSS.n12887 VSS.n12885 1.777
R16363 VSS.n12897 VSS.n12892 1.777
R16364 VSS.n12909 VSS.n12904 1.777
R16365 VSS.n12911 VSS.n12909 1.777
R16366 VSS.n12921 VSS.n12916 1.777
R16367 VSS.n12923 VSS.n12921 1.777
R16368 VSS.n12978 VSS.n12928 1.777
R16369 VSS.n12980 VSS.n12978 1.777
R16370 VSS.n12657 VSS.n12652 1.777
R16371 VSS.n12659 VSS.n12657 1.777
R16372 VSS.n12669 VSS.n12664 1.777
R16373 VSS.n12671 VSS.n12669 1.777
R16374 VSS.n12681 VSS.n12676 1.777
R16375 VSS.n12683 VSS.n12681 1.777
R16376 VSS.n12693 VSS.n12688 1.777
R16377 VSS.n12695 VSS.n12693 1.777
R16378 VSS.n12705 VSS.n12700 1.777
R16379 VSS.n12707 VSS.n12705 1.777
R16380 VSS.n12717 VSS.n12712 1.777
R16381 VSS.n12729 VSS.n12724 1.777
R16382 VSS.n12731 VSS.n12729 1.777
R16383 VSS.n12741 VSS.n12736 1.777
R16384 VSS.n12743 VSS.n12741 1.777
R16385 VSS.n12798 VSS.n12748 1.777
R16386 VSS.n12800 VSS.n12798 1.777
R16387 VSS.n9369 VSS.n9319 1.777
R16388 VSS.n9371 VSS.n9369 1.777
R16389 VSS.n9312 VSS.n9307 1.777
R16390 VSS.n9314 VSS.n9312 1.777
R16391 VSS.n9300 VSS.n9295 1.777
R16392 VSS.n9302 VSS.n9300 1.777
R16393 VSS.n9288 VSS.n9283 1.777
R16394 VSS.n9290 VSS.n9288 1.777
R16395 VSS.n9276 VSS.n9271 1.777
R16396 VSS.n9278 VSS.n9276 1.777
R16397 VSS.n9267 VSS.n9260 1.777
R16398 VSS.n9252 VSS.n9247 1.777
R16399 VSS.n9254 VSS.n9252 1.777
R16400 VSS.n9240 VSS.n9235 1.777
R16401 VSS.n9242 VSS.n9240 1.777
R16402 VSS.n9228 VSS.n9223 1.777
R16403 VSS.n9230 VSS.n9228 1.777
R16404 VSS.n9537 VSS.n9487 1.777
R16405 VSS.n9539 VSS.n9537 1.777
R16406 VSS.n9480 VSS.n9475 1.777
R16407 VSS.n9482 VSS.n9480 1.777
R16408 VSS.n9468 VSS.n9463 1.777
R16409 VSS.n9470 VSS.n9468 1.777
R16410 VSS.n9456 VSS.n9451 1.777
R16411 VSS.n9458 VSS.n9456 1.777
R16412 VSS.n9444 VSS.n9439 1.777
R16413 VSS.n9446 VSS.n9444 1.777
R16414 VSS.n9435 VSS.n9428 1.777
R16415 VSS.n9420 VSS.n9415 1.777
R16416 VSS.n9422 VSS.n9420 1.777
R16417 VSS.n9408 VSS.n9403 1.777
R16418 VSS.n9410 VSS.n9408 1.777
R16419 VSS.n9396 VSS.n9391 1.777
R16420 VSS.n9398 VSS.n9396 1.777
R16421 VSS.n9705 VSS.n9655 1.777
R16422 VSS.n9707 VSS.n9705 1.777
R16423 VSS.n9648 VSS.n9643 1.777
R16424 VSS.n9650 VSS.n9648 1.777
R16425 VSS.n9636 VSS.n9631 1.777
R16426 VSS.n9638 VSS.n9636 1.777
R16427 VSS.n9624 VSS.n9619 1.777
R16428 VSS.n9626 VSS.n9624 1.777
R16429 VSS.n9612 VSS.n9607 1.777
R16430 VSS.n9614 VSS.n9612 1.777
R16431 VSS.n9603 VSS.n9596 1.777
R16432 VSS.n9588 VSS.n9583 1.777
R16433 VSS.n9590 VSS.n9588 1.777
R16434 VSS.n9576 VSS.n9571 1.777
R16435 VSS.n9578 VSS.n9576 1.777
R16436 VSS.n9564 VSS.n9559 1.777
R16437 VSS.n9566 VSS.n9564 1.777
R16438 VSS.n9873 VSS.n9823 1.777
R16439 VSS.n9875 VSS.n9873 1.777
R16440 VSS.n9816 VSS.n9811 1.777
R16441 VSS.n9818 VSS.n9816 1.777
R16442 VSS.n9804 VSS.n9799 1.777
R16443 VSS.n9806 VSS.n9804 1.777
R16444 VSS.n9792 VSS.n9787 1.777
R16445 VSS.n9794 VSS.n9792 1.777
R16446 VSS.n9780 VSS.n9775 1.777
R16447 VSS.n9782 VSS.n9780 1.777
R16448 VSS.n9771 VSS.n9764 1.777
R16449 VSS.n9756 VSS.n9751 1.777
R16450 VSS.n9758 VSS.n9756 1.777
R16451 VSS.n9744 VSS.n9739 1.777
R16452 VSS.n9746 VSS.n9744 1.777
R16453 VSS.n9732 VSS.n9727 1.777
R16454 VSS.n9734 VSS.n9732 1.777
R16455 VSS.n10041 VSS.n9991 1.777
R16456 VSS.n10043 VSS.n10041 1.777
R16457 VSS.n9984 VSS.n9979 1.777
R16458 VSS.n9986 VSS.n9984 1.777
R16459 VSS.n9972 VSS.n9967 1.777
R16460 VSS.n9974 VSS.n9972 1.777
R16461 VSS.n9960 VSS.n9955 1.777
R16462 VSS.n9962 VSS.n9960 1.777
R16463 VSS.n9948 VSS.n9943 1.777
R16464 VSS.n9950 VSS.n9948 1.777
R16465 VSS.n9939 VSS.n9932 1.777
R16466 VSS.n9924 VSS.n9919 1.777
R16467 VSS.n9926 VSS.n9924 1.777
R16468 VSS.n9912 VSS.n9907 1.777
R16469 VSS.n9914 VSS.n9912 1.777
R16470 VSS.n9900 VSS.n9895 1.777
R16471 VSS.n9902 VSS.n9900 1.777
R16472 VSS.n10209 VSS.n10159 1.777
R16473 VSS.n10211 VSS.n10209 1.777
R16474 VSS.n10152 VSS.n10147 1.777
R16475 VSS.n10154 VSS.n10152 1.777
R16476 VSS.n10140 VSS.n10135 1.777
R16477 VSS.n10142 VSS.n10140 1.777
R16478 VSS.n10128 VSS.n10123 1.777
R16479 VSS.n10130 VSS.n10128 1.777
R16480 VSS.n10116 VSS.n10111 1.777
R16481 VSS.n10118 VSS.n10116 1.777
R16482 VSS.n10107 VSS.n10100 1.777
R16483 VSS.n10092 VSS.n10087 1.777
R16484 VSS.n10094 VSS.n10092 1.777
R16485 VSS.n10080 VSS.n10075 1.777
R16486 VSS.n10082 VSS.n10080 1.777
R16487 VSS.n10068 VSS.n10063 1.777
R16488 VSS.n10070 VSS.n10068 1.777
R16489 VSS.n10377 VSS.n10327 1.777
R16490 VSS.n10379 VSS.n10377 1.777
R16491 VSS.n10320 VSS.n10315 1.777
R16492 VSS.n10322 VSS.n10320 1.777
R16493 VSS.n10308 VSS.n10303 1.777
R16494 VSS.n10310 VSS.n10308 1.777
R16495 VSS.n10296 VSS.n10291 1.777
R16496 VSS.n10298 VSS.n10296 1.777
R16497 VSS.n10284 VSS.n10279 1.777
R16498 VSS.n10286 VSS.n10284 1.777
R16499 VSS.n10275 VSS.n10268 1.777
R16500 VSS.n10260 VSS.n10255 1.777
R16501 VSS.n10262 VSS.n10260 1.777
R16502 VSS.n10248 VSS.n10243 1.777
R16503 VSS.n10250 VSS.n10248 1.777
R16504 VSS.n10236 VSS.n10231 1.777
R16505 VSS.n10238 VSS.n10236 1.777
R16506 VSS.n10545 VSS.n10494 1.777
R16507 VSS.n10547 VSS.n10545 1.777
R16508 VSS.n10487 VSS.n10482 1.777
R16509 VSS.n10489 VSS.n10487 1.777
R16510 VSS.n10475 VSS.n10470 1.777
R16511 VSS.n10477 VSS.n10475 1.777
R16512 VSS.n10463 VSS.n10458 1.777
R16513 VSS.n10465 VSS.n10463 1.777
R16514 VSS.n10451 VSS.n10446 1.777
R16515 VSS.n10453 VSS.n10451 1.777
R16516 VSS.n10442 VSS.n10435 1.777
R16517 VSS.n10427 VSS.n10422 1.777
R16518 VSS.n10429 VSS.n10427 1.777
R16519 VSS.n10415 VSS.n10410 1.777
R16520 VSS.n10417 VSS.n10415 1.777
R16521 VSS.n10403 VSS.n10398 1.777
R16522 VSS.n10405 VSS.n10403 1.777
R16523 VSS.n2379 VSS.n2378 1.777
R16524 VSS.n2380 VSS.n2379 1.777
R16525 VSS.n2454 VSS.n2453 1.777
R16526 VSS.n2453 VSS.n2325 1.777
R16527 VSS.n2445 VSS.n2444 1.777
R16528 VSS.n2444 VSS.n2442 1.777
R16529 VSS.n2438 VSS.n2388 1.777
R16530 VSS.n2438 VSS.n2436 1.777
R16531 VSS.n2432 VSS.n2392 1.777
R16532 VSS.n2432 VSS.n2430 1.777
R16533 VSS.n2426 VSS.n2396 1.777
R16534 VSS.n2420 VSS.n2314 1.777
R16535 VSS.n2420 VSS.n2419 1.777
R16536 VSS.n2415 VSS.n2402 1.777
R16537 VSS.n2415 VSS.n2413 1.777
R16538 VSS.n2409 VSS.n2407 1.777
R16539 VSS.n2409 VSS.n2408 1.777
R16540 VSS.n2469 VSS.n2468 1.777
R16541 VSS.n2470 VSS.n2469 1.777
R16542 VSS.n2544 VSS.n2543 1.777
R16543 VSS.n2543 VSS.n2235 1.777
R16544 VSS.n2535 VSS.n2534 1.777
R16545 VSS.n2534 VSS.n2532 1.777
R16546 VSS.n2528 VSS.n2478 1.777
R16547 VSS.n2528 VSS.n2526 1.777
R16548 VSS.n2522 VSS.n2482 1.777
R16549 VSS.n2522 VSS.n2520 1.777
R16550 VSS.n2516 VSS.n2486 1.777
R16551 VSS.n2510 VSS.n2224 1.777
R16552 VSS.n2510 VSS.n2509 1.777
R16553 VSS.n2505 VSS.n2492 1.777
R16554 VSS.n2505 VSS.n2503 1.777
R16555 VSS.n2499 VSS.n2497 1.777
R16556 VSS.n2499 VSS.n2498 1.777
R16557 VSS.n2559 VSS.n2558 1.777
R16558 VSS.n2560 VSS.n2559 1.777
R16559 VSS.n2634 VSS.n2633 1.777
R16560 VSS.n2633 VSS.n2145 1.777
R16561 VSS.n2625 VSS.n2624 1.777
R16562 VSS.n2624 VSS.n2622 1.777
R16563 VSS.n2618 VSS.n2568 1.777
R16564 VSS.n2618 VSS.n2616 1.777
R16565 VSS.n2612 VSS.n2572 1.777
R16566 VSS.n2612 VSS.n2610 1.777
R16567 VSS.n2606 VSS.n2576 1.777
R16568 VSS.n2600 VSS.n2134 1.777
R16569 VSS.n2600 VSS.n2599 1.777
R16570 VSS.n2595 VSS.n2582 1.777
R16571 VSS.n2595 VSS.n2593 1.777
R16572 VSS.n2589 VSS.n2587 1.777
R16573 VSS.n2589 VSS.n2588 1.777
R16574 VSS.n2649 VSS.n2648 1.777
R16575 VSS.n2650 VSS.n2649 1.777
R16576 VSS.n2724 VSS.n2723 1.777
R16577 VSS.n2723 VSS.n2055 1.777
R16578 VSS.n2715 VSS.n2714 1.777
R16579 VSS.n2714 VSS.n2712 1.777
R16580 VSS.n2708 VSS.n2658 1.777
R16581 VSS.n2708 VSS.n2706 1.777
R16582 VSS.n2702 VSS.n2662 1.777
R16583 VSS.n2702 VSS.n2700 1.777
R16584 VSS.n2696 VSS.n2666 1.777
R16585 VSS.n2690 VSS.n2044 1.777
R16586 VSS.n2690 VSS.n2689 1.777
R16587 VSS.n2685 VSS.n2672 1.777
R16588 VSS.n2685 VSS.n2683 1.777
R16589 VSS.n2679 VSS.n2677 1.777
R16590 VSS.n2679 VSS.n2678 1.777
R16591 VSS.n2739 VSS.n2738 1.777
R16592 VSS.n2740 VSS.n2739 1.777
R16593 VSS.n2814 VSS.n2813 1.777
R16594 VSS.n2813 VSS.n1965 1.777
R16595 VSS.n2805 VSS.n2804 1.777
R16596 VSS.n2804 VSS.n2802 1.777
R16597 VSS.n2798 VSS.n2748 1.777
R16598 VSS.n2798 VSS.n2796 1.777
R16599 VSS.n2792 VSS.n2752 1.777
R16600 VSS.n2792 VSS.n2790 1.777
R16601 VSS.n2786 VSS.n2756 1.777
R16602 VSS.n2780 VSS.n1954 1.777
R16603 VSS.n2780 VSS.n2779 1.777
R16604 VSS.n2775 VSS.n2762 1.777
R16605 VSS.n2775 VSS.n2773 1.777
R16606 VSS.n2769 VSS.n2767 1.777
R16607 VSS.n2769 VSS.n2768 1.777
R16608 VSS.n2829 VSS.n2828 1.777
R16609 VSS.n2830 VSS.n2829 1.777
R16610 VSS.n2904 VSS.n2903 1.777
R16611 VSS.n2903 VSS.n1875 1.777
R16612 VSS.n2895 VSS.n2894 1.777
R16613 VSS.n2894 VSS.n2892 1.777
R16614 VSS.n2888 VSS.n2838 1.777
R16615 VSS.n2888 VSS.n2886 1.777
R16616 VSS.n2882 VSS.n2842 1.777
R16617 VSS.n2882 VSS.n2880 1.777
R16618 VSS.n2876 VSS.n2846 1.777
R16619 VSS.n2870 VSS.n1864 1.777
R16620 VSS.n2870 VSS.n2869 1.777
R16621 VSS.n2865 VSS.n2852 1.777
R16622 VSS.n2865 VSS.n2863 1.777
R16623 VSS.n2859 VSS.n2857 1.777
R16624 VSS.n2859 VSS.n2858 1.777
R16625 VSS.n2919 VSS.n2918 1.777
R16626 VSS.n2920 VSS.n2919 1.777
R16627 VSS.n2994 VSS.n2993 1.777
R16628 VSS.n2993 VSS.n1785 1.777
R16629 VSS.n2985 VSS.n2984 1.777
R16630 VSS.n2984 VSS.n2982 1.777
R16631 VSS.n2978 VSS.n2928 1.777
R16632 VSS.n2978 VSS.n2976 1.777
R16633 VSS.n2972 VSS.n2932 1.777
R16634 VSS.n2972 VSS.n2970 1.777
R16635 VSS.n2966 VSS.n2936 1.777
R16636 VSS.n2960 VSS.n1774 1.777
R16637 VSS.n2960 VSS.n2959 1.777
R16638 VSS.n2955 VSS.n2942 1.777
R16639 VSS.n2955 VSS.n2953 1.777
R16640 VSS.n2949 VSS.n2947 1.777
R16641 VSS.n2949 VSS.n2948 1.777
R16642 VSS.n3009 VSS.n3008 1.777
R16643 VSS.n3010 VSS.n3009 1.777
R16644 VSS.n3084 VSS.n3083 1.777
R16645 VSS.n3083 VSS.n1695 1.777
R16646 VSS.n3075 VSS.n3074 1.777
R16647 VSS.n3074 VSS.n3072 1.777
R16648 VSS.n3068 VSS.n3018 1.777
R16649 VSS.n3068 VSS.n3066 1.777
R16650 VSS.n3062 VSS.n3022 1.777
R16651 VSS.n3062 VSS.n3060 1.777
R16652 VSS.n3056 VSS.n3026 1.777
R16653 VSS.n3050 VSS.n1684 1.777
R16654 VSS.n3050 VSS.n3049 1.777
R16655 VSS.n3045 VSS.n3032 1.777
R16656 VSS.n3045 VSS.n3043 1.777
R16657 VSS.n3039 VSS.n3037 1.777
R16658 VSS.n3039 VSS.n3038 1.777
R16659 VSS.n6127 VSS.n6075 1.777
R16660 VSS.n6128 VSS.n6127 1.777
R16661 VSS.n6135 VSS.n6124 1.777
R16662 VSS.n6136 VSS.n6135 1.777
R16663 VSS.n6143 VSS.n6122 1.777
R16664 VSS.n6144 VSS.n6143 1.777
R16665 VSS.n6151 VSS.n6120 1.777
R16666 VSS.n6152 VSS.n6151 1.777
R16667 VSS.n6159 VSS.n6118 1.777
R16668 VSS.n6160 VSS.n6159 1.777
R16669 VSS.n6167 VSS.n6116 1.777
R16670 VSS.n6175 VSS.n6114 1.777
R16671 VSS.n6176 VSS.n6175 1.777
R16672 VSS.n6183 VSS.n6112 1.777
R16673 VSS.n6184 VSS.n6183 1.777
R16674 VSS.n6245 VSS.n6109 1.777
R16675 VSS.n6245 VSS.n6110 1.777
R16676 VSS.n6011 VSS.n5959 1.777
R16677 VSS.n6012 VSS.n6011 1.777
R16678 VSS.n6019 VSS.n6008 1.777
R16679 VSS.n6020 VSS.n6019 1.777
R16680 VSS.n6027 VSS.n6006 1.777
R16681 VSS.n6028 VSS.n6027 1.777
R16682 VSS.n6035 VSS.n6004 1.777
R16683 VSS.n6036 VSS.n6035 1.777
R16684 VSS.n6043 VSS.n6002 1.777
R16685 VSS.n6044 VSS.n6043 1.777
R16686 VSS.n6051 VSS.n6000 1.777
R16687 VSS.n6059 VSS.n5998 1.777
R16688 VSS.n6060 VSS.n6059 1.777
R16689 VSS.n6067 VSS.n5996 1.777
R16690 VSS.n6068 VSS.n6067 1.777
R16691 VSS.n6309 VSS.n5993 1.777
R16692 VSS.n6309 VSS.n5994 1.777
R16693 VSS.n5895 VSS.n5843 1.777
R16694 VSS.n5896 VSS.n5895 1.777
R16695 VSS.n5903 VSS.n5892 1.777
R16696 VSS.n5904 VSS.n5903 1.777
R16697 VSS.n5911 VSS.n5890 1.777
R16698 VSS.n5912 VSS.n5911 1.777
R16699 VSS.n5919 VSS.n5888 1.777
R16700 VSS.n5920 VSS.n5919 1.777
R16701 VSS.n5927 VSS.n5886 1.777
R16702 VSS.n5928 VSS.n5927 1.777
R16703 VSS.n5935 VSS.n5884 1.777
R16704 VSS.n5943 VSS.n5882 1.777
R16705 VSS.n5944 VSS.n5943 1.777
R16706 VSS.n5951 VSS.n5880 1.777
R16707 VSS.n5952 VSS.n5951 1.777
R16708 VSS.n6373 VSS.n5877 1.777
R16709 VSS.n6373 VSS.n5878 1.777
R16710 VSS.n7043 VSS.n5787 1.777
R16711 VSS.n7043 VSS.n5788 1.777
R16712 VSS.n7038 VSS.n7037 1.777
R16713 VSS.n7037 VSS.n5792 1.777
R16714 VSS.n7032 VSS.n7031 1.777
R16715 VSS.n7031 VSS.n5797 1.777
R16716 VSS.n7026 VSS.n7025 1.777
R16717 VSS.n7025 VSS.n5803 1.777
R16718 VSS.n7020 VSS.n7019 1.777
R16719 VSS.n7019 VSS.n5809 1.777
R16720 VSS.n7014 VSS.n7013 1.777
R16721 VSS.n7008 VSS.n7007 1.777
R16722 VSS.n7007 VSS.n5820 1.777
R16723 VSS.n7002 VSS.n7001 1.777
R16724 VSS.n7001 VSS.n5827 1.777
R16725 VSS.n6996 VSS.n6995 1.777
R16726 VSS.n6995 VSS.n5833 1.777
R16727 VSS.n6853 VSS.n6852 1.777
R16728 VSS.n6854 VSS.n6853 1.777
R16729 VSS.n6927 VSS.n6926 1.777
R16730 VSS.n6926 VSS.n6439 1.777
R16731 VSS.n6918 VSS.n6917 1.777
R16732 VSS.n6917 VSS.n6915 1.777
R16733 VSS.n6911 VSS.n6862 1.777
R16734 VSS.n6911 VSS.n6909 1.777
R16735 VSS.n6905 VSS.n6866 1.777
R16736 VSS.n6905 VSS.n6903 1.777
R16737 VSS.n6899 VSS.n6870 1.777
R16738 VSS.n6893 VSS.n6874 1.777
R16739 VSS.n6893 VSS.n6891 1.777
R16740 VSS.n6887 VSS.n6428 1.777
R16741 VSS.n6887 VSS.n6886 1.777
R16742 VSS.n6882 VSS.n6880 1.777
R16743 VSS.n6882 VSS.n6881 1.777
R16744 VSS.n6763 VSS.n6762 1.777
R16745 VSS.n6764 VSS.n6763 1.777
R16746 VSS.n6837 VSS.n6836 1.777
R16747 VSS.n6836 VSS.n6529 1.777
R16748 VSS.n6828 VSS.n6827 1.777
R16749 VSS.n6827 VSS.n6825 1.777
R16750 VSS.n6821 VSS.n6772 1.777
R16751 VSS.n6821 VSS.n6819 1.777
R16752 VSS.n6815 VSS.n6776 1.777
R16753 VSS.n6815 VSS.n6813 1.777
R16754 VSS.n6809 VSS.n6780 1.777
R16755 VSS.n6803 VSS.n6784 1.777
R16756 VSS.n6803 VSS.n6801 1.777
R16757 VSS.n6797 VSS.n6518 1.777
R16758 VSS.n6797 VSS.n6796 1.777
R16759 VSS.n6792 VSS.n6790 1.777
R16760 VSS.n6792 VSS.n6791 1.777
R16761 VSS.n6673 VSS.n6672 1.777
R16762 VSS.n6674 VSS.n6673 1.777
R16763 VSS.n6747 VSS.n6746 1.777
R16764 VSS.n6746 VSS.n6619 1.777
R16765 VSS.n6738 VSS.n6737 1.777
R16766 VSS.n6737 VSS.n6735 1.777
R16767 VSS.n6731 VSS.n6682 1.777
R16768 VSS.n6731 VSS.n6729 1.777
R16769 VSS.n6725 VSS.n6686 1.777
R16770 VSS.n6725 VSS.n6723 1.777
R16771 VSS.n6719 VSS.n6690 1.777
R16772 VSS.n6713 VSS.n6694 1.777
R16773 VSS.n6713 VSS.n6711 1.777
R16774 VSS.n6707 VSS.n6608 1.777
R16775 VSS.n6707 VSS.n6706 1.777
R16776 VSS.n6702 VSS.n6700 1.777
R16777 VSS.n6702 VSS.n6701 1.777
R16778 VSS.n17766 VSS.n17765 1.7
R16779 VSS.n5132 VSS.n3094 1.58
R16780 VSS.n17769 VSS 1.513
R16781 VSS.n397 VSS.n365 1.505
R16782 VSS.n397 VSS.n366 1.505
R16783 VSS.n418 VSS.n354 1.505
R16784 VSS.n418 VSS.n352 1.505
R16785 VSS.n18189 VSS.n18157 1.505
R16786 VSS.n18189 VSS.n18158 1.505
R16787 VSS.n18211 VSS.n18144 1.505
R16788 VSS.n18211 VSS.n18146 1.505
R16789 VSS.n5785 VSS.n518 1.504
R16790 VSS.n18230 VSS 1.458
R16791 VSS.n17769 VSS.n17768 1.361
R16792 VSS.n473 VSS 1.319
R16793 VSS.n486 VSS 1.319
R16794 VSS.n322 VSS 1.319
R16795 VSS.n17762 VSS 1.319
R16796 VSS.n17437 VSS.n17436 1.309
R16797 VSS.n17269 VSS.n17268 1.309
R16798 VSS.n17101 VSS.n17100 1.309
R16799 VSS.n16933 VSS.n16932 1.309
R16800 VSS.n16765 VSS.n16764 1.309
R16801 VSS.n16597 VSS.n16596 1.309
R16802 VSS.n10402 VSS.n10401 1.309
R16803 VSS.n6247 VSS.n6246 1.309
R16804 VSS.n6311 VSS.n6310 1.309
R16805 VSS.n6375 VSS.n6374 1.309
R16806 VSS.n6994 VSS.n5837 1.309
R16807 VSS.n16388 VSS.n16381 1.292
R16808 VSS.n16390 VSS.n16388 1.292
R16809 VSS.n16402 VSS.n16395 1.292
R16810 VSS.n16404 VSS.n16402 1.292
R16811 VSS.n16416 VSS.n16409 1.292
R16812 VSS.n16418 VSS.n16416 1.292
R16813 VSS.n16430 VSS.n16423 1.292
R16814 VSS.n16432 VSS.n16430 1.292
R16815 VSS.n16444 VSS.n16437 1.292
R16816 VSS.n16446 VSS.n16444 1.292
R16817 VSS.n16462 VSS.n16451 1.292
R16818 VSS.n16465 VSS.n16462 1.292
R16819 VSS.n16471 VSS.n14555 1.292
R16820 VSS.n16471 VSS.n14557 1.292
R16821 VSS.n16480 VSS.n14554 1.292
R16822 VSS.n16482 VSS.n16480 1.292
R16823 VSS.n16494 VSS.n16487 1.292
R16824 VSS.n16496 VSS.n16494 1.292
R16825 VSS.n16508 VSS.n16501 1.292
R16826 VSS.n16510 VSS.n16508 1.292
R16827 VSS.n16522 VSS.n16515 1.292
R16828 VSS.n16524 VSS.n16522 1.292
R16829 VSS.n16583 VSS.n16574 1.292
R16830 VSS.n16585 VSS.n16583 1.292
R16831 VSS.n16132 VSS.n16125 1.292
R16832 VSS.n16134 VSS.n16132 1.292
R16833 VSS.n16146 VSS.n16139 1.292
R16834 VSS.n16148 VSS.n16146 1.292
R16835 VSS.n16160 VSS.n16153 1.292
R16836 VSS.n16162 VSS.n16160 1.292
R16837 VSS.n16174 VSS.n16167 1.292
R16838 VSS.n16176 VSS.n16174 1.292
R16839 VSS.n16188 VSS.n16181 1.292
R16840 VSS.n16190 VSS.n16188 1.292
R16841 VSS.n16206 VSS.n16195 1.292
R16842 VSS.n16209 VSS.n16206 1.292
R16843 VSS.n16215 VSS.n14561 1.292
R16844 VSS.n16215 VSS.n14563 1.292
R16845 VSS.n16224 VSS.n14560 1.292
R16846 VSS.n16226 VSS.n16224 1.292
R16847 VSS.n16238 VSS.n16231 1.292
R16848 VSS.n16240 VSS.n16238 1.292
R16849 VSS.n16252 VSS.n16245 1.292
R16850 VSS.n16254 VSS.n16252 1.292
R16851 VSS.n16266 VSS.n16259 1.292
R16852 VSS.n16268 VSS.n16266 1.292
R16853 VSS.n16284 VSS.n16273 1.292
R16854 VSS.n16285 VSS.n16284 1.292
R16855 VSS.n15888 VSS.n15881 1.292
R16856 VSS.n15890 VSS.n15888 1.292
R16857 VSS.n15902 VSS.n15895 1.292
R16858 VSS.n15904 VSS.n15902 1.292
R16859 VSS.n15916 VSS.n15909 1.292
R16860 VSS.n15918 VSS.n15916 1.292
R16861 VSS.n15930 VSS.n15923 1.292
R16862 VSS.n15932 VSS.n15930 1.292
R16863 VSS.n15944 VSS.n15937 1.292
R16864 VSS.n15946 VSS.n15944 1.292
R16865 VSS.n15962 VSS.n15951 1.292
R16866 VSS.n15965 VSS.n15962 1.292
R16867 VSS.n15971 VSS.n14567 1.292
R16868 VSS.n15971 VSS.n14569 1.292
R16869 VSS.n15980 VSS.n14566 1.292
R16870 VSS.n15982 VSS.n15980 1.292
R16871 VSS.n15994 VSS.n15987 1.292
R16872 VSS.n15996 VSS.n15994 1.292
R16873 VSS.n16008 VSS.n16001 1.292
R16874 VSS.n16010 VSS.n16008 1.292
R16875 VSS.n16022 VSS.n16015 1.292
R16876 VSS.n16024 VSS.n16022 1.292
R16877 VSS.n16040 VSS.n16029 1.292
R16878 VSS.n16041 VSS.n16040 1.292
R16879 VSS.n15644 VSS.n15637 1.292
R16880 VSS.n15646 VSS.n15644 1.292
R16881 VSS.n15658 VSS.n15651 1.292
R16882 VSS.n15660 VSS.n15658 1.292
R16883 VSS.n15672 VSS.n15665 1.292
R16884 VSS.n15674 VSS.n15672 1.292
R16885 VSS.n15686 VSS.n15679 1.292
R16886 VSS.n15688 VSS.n15686 1.292
R16887 VSS.n15700 VSS.n15693 1.292
R16888 VSS.n15702 VSS.n15700 1.292
R16889 VSS.n15718 VSS.n15707 1.292
R16890 VSS.n15721 VSS.n15718 1.292
R16891 VSS.n15727 VSS.n14573 1.292
R16892 VSS.n15727 VSS.n14575 1.292
R16893 VSS.n15736 VSS.n14572 1.292
R16894 VSS.n15738 VSS.n15736 1.292
R16895 VSS.n15750 VSS.n15743 1.292
R16896 VSS.n15752 VSS.n15750 1.292
R16897 VSS.n15764 VSS.n15757 1.292
R16898 VSS.n15766 VSS.n15764 1.292
R16899 VSS.n15778 VSS.n15771 1.292
R16900 VSS.n15780 VSS.n15778 1.292
R16901 VSS.n15796 VSS.n15785 1.292
R16902 VSS.n15797 VSS.n15796 1.292
R16903 VSS.n15400 VSS.n15393 1.292
R16904 VSS.n15402 VSS.n15400 1.292
R16905 VSS.n15414 VSS.n15407 1.292
R16906 VSS.n15416 VSS.n15414 1.292
R16907 VSS.n15428 VSS.n15421 1.292
R16908 VSS.n15430 VSS.n15428 1.292
R16909 VSS.n15442 VSS.n15435 1.292
R16910 VSS.n15444 VSS.n15442 1.292
R16911 VSS.n15456 VSS.n15449 1.292
R16912 VSS.n15458 VSS.n15456 1.292
R16913 VSS.n15474 VSS.n15463 1.292
R16914 VSS.n15477 VSS.n15474 1.292
R16915 VSS.n15483 VSS.n14579 1.292
R16916 VSS.n15483 VSS.n14581 1.292
R16917 VSS.n15492 VSS.n14578 1.292
R16918 VSS.n15494 VSS.n15492 1.292
R16919 VSS.n15506 VSS.n15499 1.292
R16920 VSS.n15508 VSS.n15506 1.292
R16921 VSS.n15520 VSS.n15513 1.292
R16922 VSS.n15522 VSS.n15520 1.292
R16923 VSS.n15534 VSS.n15527 1.292
R16924 VSS.n15536 VSS.n15534 1.292
R16925 VSS.n15552 VSS.n15541 1.292
R16926 VSS.n15553 VSS.n15552 1.292
R16927 VSS.n15156 VSS.n15149 1.292
R16928 VSS.n15158 VSS.n15156 1.292
R16929 VSS.n15170 VSS.n15163 1.292
R16930 VSS.n15172 VSS.n15170 1.292
R16931 VSS.n15184 VSS.n15177 1.292
R16932 VSS.n15186 VSS.n15184 1.292
R16933 VSS.n15198 VSS.n15191 1.292
R16934 VSS.n15200 VSS.n15198 1.292
R16935 VSS.n15212 VSS.n15205 1.292
R16936 VSS.n15214 VSS.n15212 1.292
R16937 VSS.n15230 VSS.n15219 1.292
R16938 VSS.n15233 VSS.n15230 1.292
R16939 VSS.n15239 VSS.n14585 1.292
R16940 VSS.n15239 VSS.n14587 1.292
R16941 VSS.n15248 VSS.n14584 1.292
R16942 VSS.n15250 VSS.n15248 1.292
R16943 VSS.n15262 VSS.n15255 1.292
R16944 VSS.n15264 VSS.n15262 1.292
R16945 VSS.n15276 VSS.n15269 1.292
R16946 VSS.n15278 VSS.n15276 1.292
R16947 VSS.n15290 VSS.n15283 1.292
R16948 VSS.n15292 VSS.n15290 1.292
R16949 VSS.n15308 VSS.n15297 1.292
R16950 VSS.n15309 VSS.n15308 1.292
R16951 VSS.n14912 VSS.n14905 1.292
R16952 VSS.n14914 VSS.n14912 1.292
R16953 VSS.n14926 VSS.n14919 1.292
R16954 VSS.n14928 VSS.n14926 1.292
R16955 VSS.n14940 VSS.n14933 1.292
R16956 VSS.n14942 VSS.n14940 1.292
R16957 VSS.n14954 VSS.n14947 1.292
R16958 VSS.n14956 VSS.n14954 1.292
R16959 VSS.n14968 VSS.n14961 1.292
R16960 VSS.n14970 VSS.n14968 1.292
R16961 VSS.n14986 VSS.n14975 1.292
R16962 VSS.n14989 VSS.n14986 1.292
R16963 VSS.n14995 VSS.n14591 1.292
R16964 VSS.n14995 VSS.n14593 1.292
R16965 VSS.n15004 VSS.n14590 1.292
R16966 VSS.n15006 VSS.n15004 1.292
R16967 VSS.n15018 VSS.n15011 1.292
R16968 VSS.n15020 VSS.n15018 1.292
R16969 VSS.n15032 VSS.n15025 1.292
R16970 VSS.n15034 VSS.n15032 1.292
R16971 VSS.n15046 VSS.n15039 1.292
R16972 VSS.n15048 VSS.n15046 1.292
R16973 VSS.n15064 VSS.n15053 1.292
R16974 VSS.n15065 VSS.n15064 1.292
R16975 VSS.n14656 VSS.n14646 1.292
R16976 VSS.n14658 VSS.n14656 1.292
R16977 VSS.n14670 VSS.n14663 1.292
R16978 VSS.n14672 VSS.n14670 1.292
R16979 VSS.n14684 VSS.n14677 1.292
R16980 VSS.n14686 VSS.n14684 1.292
R16981 VSS.n14698 VSS.n14691 1.292
R16982 VSS.n14700 VSS.n14698 1.292
R16983 VSS.n14712 VSS.n14705 1.292
R16984 VSS.n14714 VSS.n14712 1.292
R16985 VSS.n14730 VSS.n14719 1.292
R16986 VSS.n14733 VSS.n14730 1.292
R16987 VSS.n14739 VSS.n14597 1.292
R16988 VSS.n14739 VSS.n14599 1.292
R16989 VSS.n14748 VSS.n14596 1.292
R16990 VSS.n14750 VSS.n14748 1.292
R16991 VSS.n14762 VSS.n14755 1.292
R16992 VSS.n14764 VSS.n14762 1.292
R16993 VSS.n14776 VSS.n14769 1.292
R16994 VSS.n14778 VSS.n14776 1.292
R16995 VSS.n14790 VSS.n14783 1.292
R16996 VSS.n14792 VSS.n14790 1.292
R16997 VSS.n14808 VSS.n14797 1.292
R16998 VSS.n14809 VSS.n14808 1.292
R16999 VSS.n12437 VSS.n12430 1.292
R17000 VSS.n12439 VSS.n12437 1.292
R17001 VSS.n12451 VSS.n12444 1.292
R17002 VSS.n12453 VSS.n12451 1.292
R17003 VSS.n12465 VSS.n12458 1.292
R17004 VSS.n12467 VSS.n12465 1.292
R17005 VSS.n12479 VSS.n12472 1.292
R17006 VSS.n12481 VSS.n12479 1.292
R17007 VSS.n12493 VSS.n12486 1.292
R17008 VSS.n12495 VSS.n12493 1.292
R17009 VSS.n12511 VSS.n12500 1.292
R17010 VSS.n12514 VSS.n12511 1.292
R17011 VSS.n12520 VSS.n10604 1.292
R17012 VSS.n12520 VSS.n10606 1.292
R17013 VSS.n12529 VSS.n10603 1.292
R17014 VSS.n12531 VSS.n12529 1.292
R17015 VSS.n12543 VSS.n12536 1.292
R17016 VSS.n12545 VSS.n12543 1.292
R17017 VSS.n12557 VSS.n12550 1.292
R17018 VSS.n12559 VSS.n12557 1.292
R17019 VSS.n12571 VSS.n12564 1.292
R17020 VSS.n12573 VSS.n12571 1.292
R17021 VSS.n12632 VSS.n12623 1.292
R17022 VSS.n12634 VSS.n12632 1.292
R17023 VSS.n12181 VSS.n12174 1.292
R17024 VSS.n12183 VSS.n12181 1.292
R17025 VSS.n12195 VSS.n12188 1.292
R17026 VSS.n12197 VSS.n12195 1.292
R17027 VSS.n12209 VSS.n12202 1.292
R17028 VSS.n12211 VSS.n12209 1.292
R17029 VSS.n12223 VSS.n12216 1.292
R17030 VSS.n12225 VSS.n12223 1.292
R17031 VSS.n12237 VSS.n12230 1.292
R17032 VSS.n12239 VSS.n12237 1.292
R17033 VSS.n12255 VSS.n12244 1.292
R17034 VSS.n12258 VSS.n12255 1.292
R17035 VSS.n12264 VSS.n10610 1.292
R17036 VSS.n12264 VSS.n10612 1.292
R17037 VSS.n12273 VSS.n10609 1.292
R17038 VSS.n12275 VSS.n12273 1.292
R17039 VSS.n12287 VSS.n12280 1.292
R17040 VSS.n12289 VSS.n12287 1.292
R17041 VSS.n12301 VSS.n12294 1.292
R17042 VSS.n12303 VSS.n12301 1.292
R17043 VSS.n12315 VSS.n12308 1.292
R17044 VSS.n12317 VSS.n12315 1.292
R17045 VSS.n12333 VSS.n12322 1.292
R17046 VSS.n12334 VSS.n12333 1.292
R17047 VSS.n11937 VSS.n11930 1.292
R17048 VSS.n11939 VSS.n11937 1.292
R17049 VSS.n11951 VSS.n11944 1.292
R17050 VSS.n11953 VSS.n11951 1.292
R17051 VSS.n11965 VSS.n11958 1.292
R17052 VSS.n11967 VSS.n11965 1.292
R17053 VSS.n11979 VSS.n11972 1.292
R17054 VSS.n11981 VSS.n11979 1.292
R17055 VSS.n11993 VSS.n11986 1.292
R17056 VSS.n11995 VSS.n11993 1.292
R17057 VSS.n12011 VSS.n12000 1.292
R17058 VSS.n12014 VSS.n12011 1.292
R17059 VSS.n12020 VSS.n10616 1.292
R17060 VSS.n12020 VSS.n10618 1.292
R17061 VSS.n12029 VSS.n10615 1.292
R17062 VSS.n12031 VSS.n12029 1.292
R17063 VSS.n12043 VSS.n12036 1.292
R17064 VSS.n12045 VSS.n12043 1.292
R17065 VSS.n12057 VSS.n12050 1.292
R17066 VSS.n12059 VSS.n12057 1.292
R17067 VSS.n12071 VSS.n12064 1.292
R17068 VSS.n12073 VSS.n12071 1.292
R17069 VSS.n12089 VSS.n12078 1.292
R17070 VSS.n12090 VSS.n12089 1.292
R17071 VSS.n11693 VSS.n11686 1.292
R17072 VSS.n11695 VSS.n11693 1.292
R17073 VSS.n11707 VSS.n11700 1.292
R17074 VSS.n11709 VSS.n11707 1.292
R17075 VSS.n11721 VSS.n11714 1.292
R17076 VSS.n11723 VSS.n11721 1.292
R17077 VSS.n11735 VSS.n11728 1.292
R17078 VSS.n11737 VSS.n11735 1.292
R17079 VSS.n11749 VSS.n11742 1.292
R17080 VSS.n11751 VSS.n11749 1.292
R17081 VSS.n11767 VSS.n11756 1.292
R17082 VSS.n11770 VSS.n11767 1.292
R17083 VSS.n11776 VSS.n10622 1.292
R17084 VSS.n11776 VSS.n10624 1.292
R17085 VSS.n11785 VSS.n10621 1.292
R17086 VSS.n11787 VSS.n11785 1.292
R17087 VSS.n11799 VSS.n11792 1.292
R17088 VSS.n11801 VSS.n11799 1.292
R17089 VSS.n11813 VSS.n11806 1.292
R17090 VSS.n11815 VSS.n11813 1.292
R17091 VSS.n11827 VSS.n11820 1.292
R17092 VSS.n11829 VSS.n11827 1.292
R17093 VSS.n11845 VSS.n11834 1.292
R17094 VSS.n11846 VSS.n11845 1.292
R17095 VSS.n11449 VSS.n11442 1.292
R17096 VSS.n11451 VSS.n11449 1.292
R17097 VSS.n11463 VSS.n11456 1.292
R17098 VSS.n11465 VSS.n11463 1.292
R17099 VSS.n11477 VSS.n11470 1.292
R17100 VSS.n11479 VSS.n11477 1.292
R17101 VSS.n11491 VSS.n11484 1.292
R17102 VSS.n11493 VSS.n11491 1.292
R17103 VSS.n11505 VSS.n11498 1.292
R17104 VSS.n11507 VSS.n11505 1.292
R17105 VSS.n11523 VSS.n11512 1.292
R17106 VSS.n11526 VSS.n11523 1.292
R17107 VSS.n11532 VSS.n10628 1.292
R17108 VSS.n11532 VSS.n10630 1.292
R17109 VSS.n11541 VSS.n10627 1.292
R17110 VSS.n11543 VSS.n11541 1.292
R17111 VSS.n11555 VSS.n11548 1.292
R17112 VSS.n11557 VSS.n11555 1.292
R17113 VSS.n11569 VSS.n11562 1.292
R17114 VSS.n11571 VSS.n11569 1.292
R17115 VSS.n11583 VSS.n11576 1.292
R17116 VSS.n11585 VSS.n11583 1.292
R17117 VSS.n11601 VSS.n11590 1.292
R17118 VSS.n11602 VSS.n11601 1.292
R17119 VSS.n11205 VSS.n11198 1.292
R17120 VSS.n11207 VSS.n11205 1.292
R17121 VSS.n11219 VSS.n11212 1.292
R17122 VSS.n11221 VSS.n11219 1.292
R17123 VSS.n11233 VSS.n11226 1.292
R17124 VSS.n11235 VSS.n11233 1.292
R17125 VSS.n11247 VSS.n11240 1.292
R17126 VSS.n11249 VSS.n11247 1.292
R17127 VSS.n11261 VSS.n11254 1.292
R17128 VSS.n11263 VSS.n11261 1.292
R17129 VSS.n11279 VSS.n11268 1.292
R17130 VSS.n11282 VSS.n11279 1.292
R17131 VSS.n11288 VSS.n10634 1.292
R17132 VSS.n11288 VSS.n10636 1.292
R17133 VSS.n11297 VSS.n10633 1.292
R17134 VSS.n11299 VSS.n11297 1.292
R17135 VSS.n11311 VSS.n11304 1.292
R17136 VSS.n11313 VSS.n11311 1.292
R17137 VSS.n11325 VSS.n11318 1.292
R17138 VSS.n11327 VSS.n11325 1.292
R17139 VSS.n11339 VSS.n11332 1.292
R17140 VSS.n11341 VSS.n11339 1.292
R17141 VSS.n11357 VSS.n11346 1.292
R17142 VSS.n11358 VSS.n11357 1.292
R17143 VSS.n10961 VSS.n10954 1.292
R17144 VSS.n10963 VSS.n10961 1.292
R17145 VSS.n10975 VSS.n10968 1.292
R17146 VSS.n10977 VSS.n10975 1.292
R17147 VSS.n10989 VSS.n10982 1.292
R17148 VSS.n10991 VSS.n10989 1.292
R17149 VSS.n11003 VSS.n10996 1.292
R17150 VSS.n11005 VSS.n11003 1.292
R17151 VSS.n11017 VSS.n11010 1.292
R17152 VSS.n11019 VSS.n11017 1.292
R17153 VSS.n11035 VSS.n11024 1.292
R17154 VSS.n11038 VSS.n11035 1.292
R17155 VSS.n11044 VSS.n10640 1.292
R17156 VSS.n11044 VSS.n10642 1.292
R17157 VSS.n11053 VSS.n10639 1.292
R17158 VSS.n11055 VSS.n11053 1.292
R17159 VSS.n11067 VSS.n11060 1.292
R17160 VSS.n11069 VSS.n11067 1.292
R17161 VSS.n11081 VSS.n11074 1.292
R17162 VSS.n11083 VSS.n11081 1.292
R17163 VSS.n11095 VSS.n11088 1.292
R17164 VSS.n11097 VSS.n11095 1.292
R17165 VSS.n11113 VSS.n11102 1.292
R17166 VSS.n11114 VSS.n11113 1.292
R17167 VSS.n10705 VSS.n10695 1.292
R17168 VSS.n10707 VSS.n10705 1.292
R17169 VSS.n10719 VSS.n10712 1.292
R17170 VSS.n10721 VSS.n10719 1.292
R17171 VSS.n10733 VSS.n10726 1.292
R17172 VSS.n10735 VSS.n10733 1.292
R17173 VSS.n10747 VSS.n10740 1.292
R17174 VSS.n10749 VSS.n10747 1.292
R17175 VSS.n10761 VSS.n10754 1.292
R17176 VSS.n10763 VSS.n10761 1.292
R17177 VSS.n10779 VSS.n10768 1.292
R17178 VSS.n10782 VSS.n10779 1.292
R17179 VSS.n10788 VSS.n10646 1.292
R17180 VSS.n10788 VSS.n10648 1.292
R17181 VSS.n10797 VSS.n10645 1.292
R17182 VSS.n10799 VSS.n10797 1.292
R17183 VSS.n10811 VSS.n10804 1.292
R17184 VSS.n10813 VSS.n10811 1.292
R17185 VSS.n10825 VSS.n10818 1.292
R17186 VSS.n10827 VSS.n10825 1.292
R17187 VSS.n10839 VSS.n10832 1.292
R17188 VSS.n10841 VSS.n10839 1.292
R17189 VSS.n10857 VSS.n10846 1.292
R17190 VSS.n10858 VSS.n10857 1.292
R17191 VSS.n9005 VSS.n8998 1.292
R17192 VSS.n9007 VSS.n9005 1.292
R17193 VSS.n9019 VSS.n9012 1.292
R17194 VSS.n9021 VSS.n9019 1.292
R17195 VSS.n9033 VSS.n9026 1.292
R17196 VSS.n9035 VSS.n9033 1.292
R17197 VSS.n9047 VSS.n9040 1.292
R17198 VSS.n9049 VSS.n9047 1.292
R17199 VSS.n9061 VSS.n9054 1.292
R17200 VSS.n9063 VSS.n9061 1.292
R17201 VSS.n9079 VSS.n9068 1.292
R17202 VSS.n9082 VSS.n9079 1.292
R17203 VSS.n9088 VSS.n7172 1.292
R17204 VSS.n9088 VSS.n7174 1.292
R17205 VSS.n9097 VSS.n7171 1.292
R17206 VSS.n9099 VSS.n9097 1.292
R17207 VSS.n9111 VSS.n9104 1.292
R17208 VSS.n9113 VSS.n9111 1.292
R17209 VSS.n9125 VSS.n9118 1.292
R17210 VSS.n9127 VSS.n9125 1.292
R17211 VSS.n9139 VSS.n9132 1.292
R17212 VSS.n9141 VSS.n9139 1.292
R17213 VSS.n9200 VSS.n9191 1.292
R17214 VSS.n9202 VSS.n9200 1.292
R17215 VSS.n8749 VSS.n8742 1.292
R17216 VSS.n8751 VSS.n8749 1.292
R17217 VSS.n8763 VSS.n8756 1.292
R17218 VSS.n8765 VSS.n8763 1.292
R17219 VSS.n8777 VSS.n8770 1.292
R17220 VSS.n8779 VSS.n8777 1.292
R17221 VSS.n8791 VSS.n8784 1.292
R17222 VSS.n8793 VSS.n8791 1.292
R17223 VSS.n8805 VSS.n8798 1.292
R17224 VSS.n8807 VSS.n8805 1.292
R17225 VSS.n8823 VSS.n8812 1.292
R17226 VSS.n8826 VSS.n8823 1.292
R17227 VSS.n8832 VSS.n7178 1.292
R17228 VSS.n8832 VSS.n7180 1.292
R17229 VSS.n8841 VSS.n7177 1.292
R17230 VSS.n8843 VSS.n8841 1.292
R17231 VSS.n8855 VSS.n8848 1.292
R17232 VSS.n8857 VSS.n8855 1.292
R17233 VSS.n8869 VSS.n8862 1.292
R17234 VSS.n8871 VSS.n8869 1.292
R17235 VSS.n8883 VSS.n8876 1.292
R17236 VSS.n8885 VSS.n8883 1.292
R17237 VSS.n8901 VSS.n8890 1.292
R17238 VSS.n8902 VSS.n8901 1.292
R17239 VSS.n8505 VSS.n8498 1.292
R17240 VSS.n8507 VSS.n8505 1.292
R17241 VSS.n8519 VSS.n8512 1.292
R17242 VSS.n8521 VSS.n8519 1.292
R17243 VSS.n8533 VSS.n8526 1.292
R17244 VSS.n8535 VSS.n8533 1.292
R17245 VSS.n8547 VSS.n8540 1.292
R17246 VSS.n8549 VSS.n8547 1.292
R17247 VSS.n8561 VSS.n8554 1.292
R17248 VSS.n8563 VSS.n8561 1.292
R17249 VSS.n8579 VSS.n8568 1.292
R17250 VSS.n8582 VSS.n8579 1.292
R17251 VSS.n8588 VSS.n7184 1.292
R17252 VSS.n8588 VSS.n7186 1.292
R17253 VSS.n8597 VSS.n7183 1.292
R17254 VSS.n8599 VSS.n8597 1.292
R17255 VSS.n8611 VSS.n8604 1.292
R17256 VSS.n8613 VSS.n8611 1.292
R17257 VSS.n8625 VSS.n8618 1.292
R17258 VSS.n8627 VSS.n8625 1.292
R17259 VSS.n8639 VSS.n8632 1.292
R17260 VSS.n8641 VSS.n8639 1.292
R17261 VSS.n8657 VSS.n8646 1.292
R17262 VSS.n8658 VSS.n8657 1.292
R17263 VSS.n8261 VSS.n8254 1.292
R17264 VSS.n8263 VSS.n8261 1.292
R17265 VSS.n8275 VSS.n8268 1.292
R17266 VSS.n8277 VSS.n8275 1.292
R17267 VSS.n8289 VSS.n8282 1.292
R17268 VSS.n8291 VSS.n8289 1.292
R17269 VSS.n8303 VSS.n8296 1.292
R17270 VSS.n8305 VSS.n8303 1.292
R17271 VSS.n8317 VSS.n8310 1.292
R17272 VSS.n8319 VSS.n8317 1.292
R17273 VSS.n8335 VSS.n8324 1.292
R17274 VSS.n8338 VSS.n8335 1.292
R17275 VSS.n8344 VSS.n7190 1.292
R17276 VSS.n8344 VSS.n7192 1.292
R17277 VSS.n8353 VSS.n7189 1.292
R17278 VSS.n8355 VSS.n8353 1.292
R17279 VSS.n8367 VSS.n8360 1.292
R17280 VSS.n8369 VSS.n8367 1.292
R17281 VSS.n8381 VSS.n8374 1.292
R17282 VSS.n8383 VSS.n8381 1.292
R17283 VSS.n8395 VSS.n8388 1.292
R17284 VSS.n8397 VSS.n8395 1.292
R17285 VSS.n8413 VSS.n8402 1.292
R17286 VSS.n8414 VSS.n8413 1.292
R17287 VSS.n8017 VSS.n8010 1.292
R17288 VSS.n8019 VSS.n8017 1.292
R17289 VSS.n8031 VSS.n8024 1.292
R17290 VSS.n8033 VSS.n8031 1.292
R17291 VSS.n8045 VSS.n8038 1.292
R17292 VSS.n8047 VSS.n8045 1.292
R17293 VSS.n8059 VSS.n8052 1.292
R17294 VSS.n8061 VSS.n8059 1.292
R17295 VSS.n8073 VSS.n8066 1.292
R17296 VSS.n8075 VSS.n8073 1.292
R17297 VSS.n8091 VSS.n8080 1.292
R17298 VSS.n8094 VSS.n8091 1.292
R17299 VSS.n8100 VSS.n7196 1.292
R17300 VSS.n8100 VSS.n7198 1.292
R17301 VSS.n8109 VSS.n7195 1.292
R17302 VSS.n8111 VSS.n8109 1.292
R17303 VSS.n8123 VSS.n8116 1.292
R17304 VSS.n8125 VSS.n8123 1.292
R17305 VSS.n8137 VSS.n8130 1.292
R17306 VSS.n8139 VSS.n8137 1.292
R17307 VSS.n8151 VSS.n8144 1.292
R17308 VSS.n8153 VSS.n8151 1.292
R17309 VSS.n8169 VSS.n8158 1.292
R17310 VSS.n8170 VSS.n8169 1.292
R17311 VSS.n7773 VSS.n7766 1.292
R17312 VSS.n7775 VSS.n7773 1.292
R17313 VSS.n7787 VSS.n7780 1.292
R17314 VSS.n7789 VSS.n7787 1.292
R17315 VSS.n7801 VSS.n7794 1.292
R17316 VSS.n7803 VSS.n7801 1.292
R17317 VSS.n7815 VSS.n7808 1.292
R17318 VSS.n7817 VSS.n7815 1.292
R17319 VSS.n7829 VSS.n7822 1.292
R17320 VSS.n7831 VSS.n7829 1.292
R17321 VSS.n7847 VSS.n7836 1.292
R17322 VSS.n7850 VSS.n7847 1.292
R17323 VSS.n7856 VSS.n7202 1.292
R17324 VSS.n7856 VSS.n7204 1.292
R17325 VSS.n7865 VSS.n7201 1.292
R17326 VSS.n7867 VSS.n7865 1.292
R17327 VSS.n7879 VSS.n7872 1.292
R17328 VSS.n7881 VSS.n7879 1.292
R17329 VSS.n7893 VSS.n7886 1.292
R17330 VSS.n7895 VSS.n7893 1.292
R17331 VSS.n7907 VSS.n7900 1.292
R17332 VSS.n7909 VSS.n7907 1.292
R17333 VSS.n7925 VSS.n7914 1.292
R17334 VSS.n7926 VSS.n7925 1.292
R17335 VSS.n7529 VSS.n7522 1.292
R17336 VSS.n7531 VSS.n7529 1.292
R17337 VSS.n7543 VSS.n7536 1.292
R17338 VSS.n7545 VSS.n7543 1.292
R17339 VSS.n7557 VSS.n7550 1.292
R17340 VSS.n7559 VSS.n7557 1.292
R17341 VSS.n7571 VSS.n7564 1.292
R17342 VSS.n7573 VSS.n7571 1.292
R17343 VSS.n7585 VSS.n7578 1.292
R17344 VSS.n7587 VSS.n7585 1.292
R17345 VSS.n7603 VSS.n7592 1.292
R17346 VSS.n7606 VSS.n7603 1.292
R17347 VSS.n7612 VSS.n7208 1.292
R17348 VSS.n7612 VSS.n7210 1.292
R17349 VSS.n7621 VSS.n7207 1.292
R17350 VSS.n7623 VSS.n7621 1.292
R17351 VSS.n7635 VSS.n7628 1.292
R17352 VSS.n7637 VSS.n7635 1.292
R17353 VSS.n7649 VSS.n7642 1.292
R17354 VSS.n7651 VSS.n7649 1.292
R17355 VSS.n7663 VSS.n7656 1.292
R17356 VSS.n7665 VSS.n7663 1.292
R17357 VSS.n7681 VSS.n7670 1.292
R17358 VSS.n7682 VSS.n7681 1.292
R17359 VSS.n7273 VSS.n7263 1.292
R17360 VSS.n7275 VSS.n7273 1.292
R17361 VSS.n7287 VSS.n7280 1.292
R17362 VSS.n7289 VSS.n7287 1.292
R17363 VSS.n7301 VSS.n7294 1.292
R17364 VSS.n7303 VSS.n7301 1.292
R17365 VSS.n7315 VSS.n7308 1.292
R17366 VSS.n7317 VSS.n7315 1.292
R17367 VSS.n7329 VSS.n7322 1.292
R17368 VSS.n7331 VSS.n7329 1.292
R17369 VSS.n7347 VSS.n7336 1.292
R17370 VSS.n7350 VSS.n7347 1.292
R17371 VSS.n7356 VSS.n7214 1.292
R17372 VSS.n7356 VSS.n7216 1.292
R17373 VSS.n7365 VSS.n7213 1.292
R17374 VSS.n7367 VSS.n7365 1.292
R17375 VSS.n7379 VSS.n7372 1.292
R17376 VSS.n7381 VSS.n7379 1.292
R17377 VSS.n7393 VSS.n7386 1.292
R17378 VSS.n7395 VSS.n7393 1.292
R17379 VSS.n7407 VSS.n7400 1.292
R17380 VSS.n7409 VSS.n7407 1.292
R17381 VSS.n7425 VSS.n7414 1.292
R17382 VSS.n7426 VSS.n7425 1.292
R17383 VSS.n1259 VSS.n1019 1.292
R17384 VSS.n1259 VSS.n1020 1.292
R17385 VSS.n1253 VSS.n1252 1.292
R17386 VSS.n1252 VSS.n1029 1.292
R17387 VSS.n1241 VSS.n1033 1.292
R17388 VSS.n1241 VSS.n1240 1.292
R17389 VSS.n1236 VSS.n1040 1.292
R17390 VSS.n1236 VSS.n1041 1.292
R17391 VSS.n1230 VSS.n1229 1.292
R17392 VSS.n1229 VSS.n1048 1.292
R17393 VSS.n1218 VSS.n1052 1.292
R17394 VSS.n1218 VSS.n1217 1.292
R17395 VSS.n1213 VSS.n1059 1.292
R17396 VSS.n1213 VSS.n1060 1.292
R17397 VSS.n1207 VSS.n1206 1.292
R17398 VSS.n1206 VSS.n1067 1.292
R17399 VSS.n1195 VSS.n1071 1.292
R17400 VSS.n1195 VSS.n1194 1.292
R17401 VSS.n1190 VSS.n1078 1.292
R17402 VSS.n1190 VSS.n1079 1.292
R17403 VSS.n1184 VSS.n1183 1.292
R17404 VSS.n1183 VSS.n1086 1.292
R17405 VSS.n1172 VSS.n1090 1.292
R17406 VSS.n1172 VSS.n1171 1.292
R17407 VSS.n922 VSS.n921 1.292
R17408 VSS.n922 VSS.n711 1.292
R17409 VSS.n933 VSS.n706 1.292
R17410 VSS.n934 VSS.n933 1.292
R17411 VSS.n939 VSS.n938 1.292
R17412 VSS.n938 VSS.n700 1.292
R17413 VSS.n950 VSS.n696 1.292
R17414 VSS.n950 VSS.n698 1.292
R17415 VSS.n957 VSS.n956 1.292
R17416 VSS.n957 VSS.n690 1.292
R17417 VSS.n968 VSS.n685 1.292
R17418 VSS.n969 VSS.n968 1.292
R17419 VSS.n974 VSS.n973 1.292
R17420 VSS.n973 VSS.n679 1.292
R17421 VSS.n985 VSS.n675 1.292
R17422 VSS.n985 VSS.n677 1.292
R17423 VSS.n992 VSS.n991 1.292
R17424 VSS.n992 VSS.n669 1.292
R17425 VSS.n1003 VSS.n664 1.292
R17426 VSS.n1004 VSS.n1003 1.292
R17427 VSS.n1009 VSS.n1008 1.292
R17428 VSS.n1008 VSS.n658 1.292
R17429 VSS.n1266 VSS.n655 1.292
R17430 VSS.n1266 VSS.n656 1.292
R17431 VSS.n786 VSS.n778 1.292
R17432 VSS.n787 VSS.n786 1.292
R17433 VSS.n792 VSS.n791 1.292
R17434 VSS.n791 VSS.n772 1.292
R17435 VSS.n803 VSS.n768 1.292
R17436 VSS.n803 VSS.n770 1.292
R17437 VSS.n810 VSS.n809 1.292
R17438 VSS.n810 VSS.n762 1.292
R17439 VSS.n821 VSS.n757 1.292
R17440 VSS.n822 VSS.n821 1.292
R17441 VSS.n827 VSS.n826 1.292
R17442 VSS.n826 VSS.n751 1.292
R17443 VSS.n838 VSS.n747 1.292
R17444 VSS.n838 VSS.n749 1.292
R17445 VSS.n845 VSS.n844 1.292
R17446 VSS.n845 VSS.n741 1.292
R17447 VSS.n856 VSS.n736 1.292
R17448 VSS.n857 VSS.n856 1.292
R17449 VSS.n862 VSS.n861 1.292
R17450 VSS.n861 VSS.n730 1.292
R17451 VSS.n873 VSS.n725 1.292
R17452 VSS.n873 VSS.n728 1.292
R17453 VSS.n880 VSS.n721 1.292
R17454 VSS.n880 VSS.n719 1.292
R17455 VSS.n5605 VSS.n5604 1.292
R17456 VSS.n5604 VSS.n5601 1.292
R17457 VSS.n5782 VSS.n521 1.292
R17458 VSS.n5782 VSS.n522 1.292
R17459 VSS.n5776 VSS.n5775 1.292
R17460 VSS.n5775 VSS.n529 1.292
R17461 VSS.n5764 VSS.n533 1.292
R17462 VSS.n5764 VSS.n5763 1.292
R17463 VSS.n5759 VSS.n540 1.292
R17464 VSS.n5759 VSS.n541 1.292
R17465 VSS.n5753 VSS.n5752 1.292
R17466 VSS.n5752 VSS.n548 1.292
R17467 VSS.n5741 VSS.n552 1.292
R17468 VSS.n5741 VSS.n5740 1.292
R17469 VSS.n5736 VSS.n559 1.292
R17470 VSS.n5736 VSS.n560 1.292
R17471 VSS.n5730 VSS.n5729 1.292
R17472 VSS.n5729 VSS.n567 1.292
R17473 VSS.n5718 VSS.n571 1.292
R17474 VSS.n5718 VSS.n5717 1.292
R17475 VSS.n5713 VSS.n578 1.292
R17476 VSS.n5713 VSS.n579 1.292
R17477 VSS.n5707 VSS.n5706 1.292
R17478 VSS.n5706 VSS.n586 1.292
R17479 VSS.n5500 VSS.n1441 1.292
R17480 VSS.n5501 VSS.n5500 1.292
R17481 VSS.n5506 VSS.n5505 1.292
R17482 VSS.n5505 VSS.n1435 1.292
R17483 VSS.n5517 VSS.n1431 1.292
R17484 VSS.n5517 VSS.n1433 1.292
R17485 VSS.n5524 VSS.n5523 1.292
R17486 VSS.n5524 VSS.n1425 1.292
R17487 VSS.n5535 VSS.n1420 1.292
R17488 VSS.n5536 VSS.n5535 1.292
R17489 VSS.n5541 VSS.n5540 1.292
R17490 VSS.n5540 VSS.n1414 1.292
R17491 VSS.n5552 VSS.n1410 1.292
R17492 VSS.n5552 VSS.n1412 1.292
R17493 VSS.n5559 VSS.n5558 1.292
R17494 VSS.n5559 VSS.n1404 1.292
R17495 VSS.n5570 VSS.n1399 1.292
R17496 VSS.n5571 VSS.n5570 1.292
R17497 VSS.n5576 VSS.n5575 1.292
R17498 VSS.n5575 VSS.n1391 1.292
R17499 VSS.n1392 VSS.n1389 1.292
R17500 VSS.n5588 VSS.n1389 1.292
R17501 VSS.n5612 VSS.n1384 1.292
R17502 VSS.n5612 VSS.n1382 1.292
R17503 VSS.n5397 VSS.n5396 1.292
R17504 VSS.n5396 VSS.n5237 1.292
R17505 VSS.n5385 VSS.n5239 1.292
R17506 VSS.n5385 VSS.n5384 1.292
R17507 VSS.n5380 VSS.n5247 1.292
R17508 VSS.n5380 VSS.n5248 1.292
R17509 VSS.n5374 VSS.n5373 1.292
R17510 VSS.n5373 VSS.n5255 1.292
R17511 VSS.n5362 VSS.n5259 1.292
R17512 VSS.n5362 VSS.n5361 1.292
R17513 VSS.n5357 VSS.n5266 1.292
R17514 VSS.n5357 VSS.n5267 1.292
R17515 VSS.n5351 VSS.n5350 1.292
R17516 VSS.n5350 VSS.n5274 1.292
R17517 VSS.n5339 VSS.n5278 1.292
R17518 VSS.n5339 VSS.n5338 1.292
R17519 VSS.n5334 VSS.n5285 1.292
R17520 VSS.n5334 VSS.n5286 1.292
R17521 VSS.n5328 VSS.n5327 1.292
R17522 VSS.n5327 VSS.n5293 1.292
R17523 VSS.n5316 VSS.n5297 1.292
R17524 VSS.n5316 VSS.n5315 1.292
R17525 VSS.n5311 VSS.n5305 1.292
R17526 VSS.n5311 VSS.n5306 1.292
R17527 VSS.n5141 VSS.n1582 1.292
R17528 VSS.n5142 VSS.n5141 1.292
R17529 VSS.n5147 VSS.n5146 1.292
R17530 VSS.n5146 VSS.n1576 1.292
R17531 VSS.n5158 VSS.n1572 1.292
R17532 VSS.n5158 VSS.n1574 1.292
R17533 VSS.n5165 VSS.n5164 1.292
R17534 VSS.n5165 VSS.n1566 1.292
R17535 VSS.n5176 VSS.n1561 1.292
R17536 VSS.n5177 VSS.n5176 1.292
R17537 VSS.n5182 VSS.n5181 1.292
R17538 VSS.n5181 VSS.n1555 1.292
R17539 VSS.n5193 VSS.n1551 1.292
R17540 VSS.n5193 VSS.n1553 1.292
R17541 VSS.n5200 VSS.n5199 1.292
R17542 VSS.n5200 VSS.n1545 1.292
R17543 VSS.n5211 VSS.n1540 1.292
R17544 VSS.n5212 VSS.n5211 1.292
R17545 VSS.n5217 VSS.n5216 1.292
R17546 VSS.n5216 VSS.n1532 1.292
R17547 VSS.n1533 VSS.n1530 1.292
R17548 VSS.n5229 VSS.n1530 1.292
R17549 VSS.n5404 VSS.n1525 1.292
R17550 VSS.n5404 VSS.n1523 1.292
R17551 VSS.n4926 VSS.n4762 1.292
R17552 VSS.n4926 VSS.n4763 1.292
R17553 VSS.n4920 VSS.n4919 1.292
R17554 VSS.n4919 VSS.n4773 1.292
R17555 VSS.n4908 VSS.n4777 1.292
R17556 VSS.n4908 VSS.n4907 1.292
R17557 VSS.n4903 VSS.n4784 1.292
R17558 VSS.n4903 VSS.n4785 1.292
R17559 VSS.n4897 VSS.n4896 1.292
R17560 VSS.n4896 VSS.n4792 1.292
R17561 VSS.n4885 VSS.n4796 1.292
R17562 VSS.n4885 VSS.n4884 1.292
R17563 VSS.n4880 VSS.n4803 1.292
R17564 VSS.n4880 VSS.n4804 1.292
R17565 VSS.n4874 VSS.n4873 1.292
R17566 VSS.n4873 VSS.n4811 1.292
R17567 VSS.n4862 VSS.n4815 1.292
R17568 VSS.n4862 VSS.n4861 1.292
R17569 VSS.n4857 VSS.n4822 1.292
R17570 VSS.n4857 VSS.n4823 1.292
R17571 VSS.n4851 VSS.n4850 1.292
R17572 VSS.n4850 VSS.n4830 1.292
R17573 VSS.n4839 VSS.n4834 1.292
R17574 VSS.n4839 VSS.n4838 1.292
R17575 VSS.n5019 VSS.n4651 1.292
R17576 VSS.n5019 VSS.n4652 1.292
R17577 VSS.n5013 VSS.n5012 1.292
R17578 VSS.n5012 VSS.n4661 1.292
R17579 VSS.n5001 VSS.n4665 1.292
R17580 VSS.n5001 VSS.n5000 1.292
R17581 VSS.n4996 VSS.n4672 1.292
R17582 VSS.n4996 VSS.n4673 1.292
R17583 VSS.n4990 VSS.n4989 1.292
R17584 VSS.n4989 VSS.n4680 1.292
R17585 VSS.n4978 VSS.n4684 1.292
R17586 VSS.n4978 VSS.n4977 1.292
R17587 VSS.n4973 VSS.n4691 1.292
R17588 VSS.n4973 VSS.n4692 1.292
R17589 VSS.n4967 VSS.n4966 1.292
R17590 VSS.n4966 VSS.n4699 1.292
R17591 VSS.n4955 VSS.n4703 1.292
R17592 VSS.n4955 VSS.n4954 1.292
R17593 VSS.n4950 VSS.n4710 1.292
R17594 VSS.n4950 VSS.n4711 1.292
R17595 VSS.n4944 VSS.n4943 1.292
R17596 VSS.n4943 VSS.n4718 1.292
R17597 VSS.n4932 VSS.n4722 1.292
R17598 VSS.n4932 VSS.n4931 1.292
R17599 VSS.n4547 VSS.n4546 1.292
R17600 VSS.n4546 VSS.n3214 1.292
R17601 VSS.n4558 VSS.n3210 1.292
R17602 VSS.n4558 VSS.n3212 1.292
R17603 VSS.n4565 VSS.n4564 1.292
R17604 VSS.n4565 VSS.n3204 1.292
R17605 VSS.n4576 VSS.n3199 1.292
R17606 VSS.n4577 VSS.n4576 1.292
R17607 VSS.n4582 VSS.n4581 1.292
R17608 VSS.n4581 VSS.n3193 1.292
R17609 VSS.n4593 VSS.n3189 1.292
R17610 VSS.n4593 VSS.n3191 1.292
R17611 VSS.n4600 VSS.n4599 1.292
R17612 VSS.n4600 VSS.n3183 1.292
R17613 VSS.n4611 VSS.n3178 1.292
R17614 VSS.n4612 VSS.n4611 1.292
R17615 VSS.n4617 VSS.n4616 1.292
R17616 VSS.n4616 VSS.n3172 1.292
R17617 VSS.n4628 VSS.n3168 1.292
R17618 VSS.n4628 VSS.n3170 1.292
R17619 VSS.n4635 VSS.n4634 1.292
R17620 VSS.n4635 VSS.n3162 1.292
R17621 VSS.n4646 VSS.n3158 1.292
R17622 VSS.n4647 VSS.n4646 1.292
R17623 VSS.n4317 VSS.n4172 1.292
R17624 VSS.n4317 VSS.n4173 1.292
R17625 VSS.n4311 VSS.n4310 1.292
R17626 VSS.n4310 VSS.n4183 1.292
R17627 VSS.n4299 VSS.n4187 1.292
R17628 VSS.n4299 VSS.n4298 1.292
R17629 VSS.n4294 VSS.n4194 1.292
R17630 VSS.n4294 VSS.n4195 1.292
R17631 VSS.n4288 VSS.n4287 1.292
R17632 VSS.n4287 VSS.n4202 1.292
R17633 VSS.n4276 VSS.n4206 1.292
R17634 VSS.n4276 VSS.n4275 1.292
R17635 VSS.n4271 VSS.n4213 1.292
R17636 VSS.n4271 VSS.n4214 1.292
R17637 VSS.n4265 VSS.n4264 1.292
R17638 VSS.n4264 VSS.n4221 1.292
R17639 VSS.n4253 VSS.n4225 1.292
R17640 VSS.n4253 VSS.n4252 1.292
R17641 VSS.n4248 VSS.n4232 1.292
R17642 VSS.n4248 VSS.n4233 1.292
R17643 VSS.n4242 VSS.n4241 1.292
R17644 VSS.n4241 VSS.n3223 1.292
R17645 VSS.n3224 VSS.n3221 1.292
R17646 VSS.n4541 VSS.n3221 1.292
R17647 VSS.n4410 VSS.n4061 1.292
R17648 VSS.n4410 VSS.n4062 1.292
R17649 VSS.n4404 VSS.n4403 1.292
R17650 VSS.n4403 VSS.n4071 1.292
R17651 VSS.n4392 VSS.n4075 1.292
R17652 VSS.n4392 VSS.n4391 1.292
R17653 VSS.n4387 VSS.n4082 1.292
R17654 VSS.n4387 VSS.n4083 1.292
R17655 VSS.n4381 VSS.n4380 1.292
R17656 VSS.n4380 VSS.n4090 1.292
R17657 VSS.n4369 VSS.n4094 1.292
R17658 VSS.n4369 VSS.n4368 1.292
R17659 VSS.n4364 VSS.n4101 1.292
R17660 VSS.n4364 VSS.n4102 1.292
R17661 VSS.n4358 VSS.n4357 1.292
R17662 VSS.n4357 VSS.n4109 1.292
R17663 VSS.n4346 VSS.n4113 1.292
R17664 VSS.n4346 VSS.n4345 1.292
R17665 VSS.n4341 VSS.n4120 1.292
R17666 VSS.n4341 VSS.n4121 1.292
R17667 VSS.n4335 VSS.n4334 1.292
R17668 VSS.n4334 VSS.n4128 1.292
R17669 VSS.n4323 VSS.n4132 1.292
R17670 VSS.n4323 VSS.n4322 1.292
R17671 VSS.n3964 VSS.n3963 1.292
R17672 VSS.n3964 VSS.n3381 1.292
R17673 VSS.n3975 VSS.n3376 1.292
R17674 VSS.n3976 VSS.n3975 1.292
R17675 VSS.n3981 VSS.n3980 1.292
R17676 VSS.n3980 VSS.n3370 1.292
R17677 VSS.n3992 VSS.n3366 1.292
R17678 VSS.n3992 VSS.n3368 1.292
R17679 VSS.n3999 VSS.n3998 1.292
R17680 VSS.n3999 VSS.n3360 1.292
R17681 VSS.n4010 VSS.n3355 1.292
R17682 VSS.n4011 VSS.n4010 1.292
R17683 VSS.n4016 VSS.n4015 1.292
R17684 VSS.n4015 VSS.n3349 1.292
R17685 VSS.n4027 VSS.n3345 1.292
R17686 VSS.n4027 VSS.n3347 1.292
R17687 VSS.n4034 VSS.n4033 1.292
R17688 VSS.n4034 VSS.n3339 1.292
R17689 VSS.n4045 VSS.n3334 1.292
R17690 VSS.n4046 VSS.n4045 1.292
R17691 VSS.n4051 VSS.n4050 1.292
R17692 VSS.n4050 VSS.n3328 1.292
R17693 VSS.n4417 VSS.n3325 1.292
R17694 VSS.n4417 VSS.n3326 1.292
R17695 VSS.n3713 VSS.n3560 1.292
R17696 VSS.n3713 VSS.n3561 1.292
R17697 VSS.n3707 VSS.n3706 1.292
R17698 VSS.n3706 VSS.n3571 1.292
R17699 VSS.n3695 VSS.n3575 1.292
R17700 VSS.n3695 VSS.n3694 1.292
R17701 VSS.n3690 VSS.n3582 1.292
R17702 VSS.n3690 VSS.n3583 1.292
R17703 VSS.n3684 VSS.n3683 1.292
R17704 VSS.n3683 VSS.n3590 1.292
R17705 VSS.n3672 VSS.n3594 1.292
R17706 VSS.n3672 VSS.n3671 1.292
R17707 VSS.n3667 VSS.n3601 1.292
R17708 VSS.n3667 VSS.n3602 1.292
R17709 VSS.n3661 VSS.n3660 1.292
R17710 VSS.n3660 VSS.n3609 1.292
R17711 VSS.n3649 VSS.n3613 1.292
R17712 VSS.n3649 VSS.n3648 1.292
R17713 VSS.n3644 VSS.n3620 1.292
R17714 VSS.n3644 VSS.n3621 1.292
R17715 VSS.n3638 VSS.n3637 1.292
R17716 VSS.n3637 VSS.n3632 1.292
R17717 VSS.n3956 VSS.n3389 1.292
R17718 VSS.n3956 VSS.n3390 1.292
R17719 VSS.n3807 VSS.n3806 1.292
R17720 VSS.n3806 VSS.n3452 1.292
R17721 VSS.n3800 VSS.n3799 1.292
R17722 VSS.n3799 VSS.n3458 1.292
R17723 VSS.n3788 VSS.n3463 1.292
R17724 VSS.n3788 VSS.n3787 1.292
R17725 VSS.n3783 VSS.n3470 1.292
R17726 VSS.n3783 VSS.n3471 1.292
R17727 VSS.n3777 VSS.n3776 1.292
R17728 VSS.n3776 VSS.n3478 1.292
R17729 VSS.n3765 VSS.n3482 1.292
R17730 VSS.n3765 VSS.n3764 1.292
R17731 VSS.n3760 VSS.n3489 1.292
R17732 VSS.n3760 VSS.n3490 1.292
R17733 VSS.n3754 VSS.n3753 1.292
R17734 VSS.n3753 VSS.n3497 1.292
R17735 VSS.n3742 VSS.n3501 1.292
R17736 VSS.n3742 VSS.n3741 1.292
R17737 VSS.n3737 VSS.n3508 1.292
R17738 VSS.n3737 VSS.n3509 1.292
R17739 VSS.n3731 VSS.n3730 1.292
R17740 VSS.n3730 VSS.n3516 1.292
R17741 VSS.n3719 VSS.n3520 1.292
R17742 VSS.n3719 VSS.n3718 1.292
R17743 VSS.n17866 VSS 1.292
R17744 VSS.n17753 VSS 1.283
R17745 VSS.n16377 VSS.n16375 1.28
R17746 VSS.n16121 VSS.n16120 1.28
R17747 VSS.n15877 VSS.n15875 1.28
R17748 VSS.n15633 VSS.n15632 1.28
R17749 VSS.n15389 VSS.n15387 1.28
R17750 VSS.n15145 VSS.n15144 1.28
R17751 VSS.n14901 VSS.n14899 1.28
R17752 VSS.n12426 VSS.n12424 1.28
R17753 VSS.n12170 VSS.n12169 1.28
R17754 VSS.n11926 VSS.n11924 1.28
R17755 VSS.n11682 VSS.n11681 1.28
R17756 VSS.n11438 VSS.n11436 1.28
R17757 VSS.n11194 VSS.n11193 1.28
R17758 VSS.n10950 VSS.n10948 1.28
R17759 VSS.n8994 VSS.n8992 1.28
R17760 VSS.n8738 VSS.n8737 1.28
R17761 VSS.n8494 VSS.n8492 1.28
R17762 VSS.n8250 VSS.n8249 1.28
R17763 VSS.n8006 VSS.n8004 1.28
R17764 VSS.n7762 VSS.n7761 1.28
R17765 VSS.n7518 VSS.n7516 1.28
R17766 VSS.n1272 VSS.n650 1.28
R17767 VSS.n914 VSS.n885 1.28
R17768 VSS.n5701 VSS.n5700 1.28
R17769 VSS.n5618 VSS.n5617 1.28
R17770 VSS.n5493 VSS.n5492 1.28
R17771 VSS.n5410 VSS.n5409 1.28
R17772 VSS.n4760 VSS.n4759 1.28
R17773 VSS.n5023 VSS.n5022 1.28
R17774 VSS.n4543 VSS.n3220 1.28
R17775 VSS.n4170 VSS.n4169 1.28
R17776 VSS.n4423 VSS.n3320 1.28
R17777 VSS.n3951 VSS.n3950 1.28
R17778 VSS.n3558 VSS.n3557 1.28
R17779 VSS.n14315 VSS.n14314 1.244
R17780 VSS.n14322 VSS.n14321 1.244
R17781 VSS.n14327 VSS.n14326 1.244
R17782 VSS.n14334 VSS.n14333 1.244
R17783 VSS.n14339 VSS.n14338 1.244
R17784 VSS.n14346 VSS.n14345 1.244
R17785 VSS.n14351 VSS.n14350 1.244
R17786 VSS.n14358 VSS.n14357 1.244
R17787 VSS.n14363 VSS.n14362 1.244
R17788 VSS.n14370 VSS.n14369 1.244
R17789 VSS.n14375 VSS.n14374 1.244
R17790 VSS VSS.n14380 1.244
R17791 VSS.n14382 VSS.n14381 1.244
R17792 VSS.n14387 VSS.n14386 1.244
R17793 VSS.n14394 VSS.n14393 1.244
R17794 VSS.n14399 VSS.n14398 1.244
R17795 VSS.n14406 VSS.n14405 1.244
R17796 VSS.n14411 VSS.n14410 1.244
R17797 VSS.n14463 VSS.n14462 1.244
R17798 VSS.n14135 VSS.n14134 1.244
R17799 VSS.n14142 VSS.n14141 1.244
R17800 VSS.n14147 VSS.n14146 1.244
R17801 VSS.n14154 VSS.n14153 1.244
R17802 VSS.n14159 VSS.n14158 1.244
R17803 VSS.n14166 VSS.n14165 1.244
R17804 VSS.n14171 VSS.n14170 1.244
R17805 VSS.n14178 VSS.n14177 1.244
R17806 VSS.n14183 VSS.n14182 1.244
R17807 VSS.n14190 VSS.n14189 1.244
R17808 VSS.n14195 VSS.n14194 1.244
R17809 VSS VSS.n14200 1.244
R17810 VSS.n14202 VSS.n14201 1.244
R17811 VSS.n14207 VSS.n14206 1.244
R17812 VSS.n14214 VSS.n14213 1.244
R17813 VSS.n14219 VSS.n14218 1.244
R17814 VSS.n14226 VSS.n14225 1.244
R17815 VSS.n14231 VSS.n14230 1.244
R17816 VSS.n14283 VSS.n14282 1.244
R17817 VSS.n17529 VSS.n17528 1.244
R17818 VSS.n17583 VSS.n17582 1.244
R17819 VSS.n17517 VSS.n17516 1.244
R17820 VSS.n17524 VSS.n17523 1.244
R17821 VSS.n17505 VSS.n17504 1.244
R17822 VSS.n17512 VSS.n17511 1.244
R17823 VSS.n17493 VSS.n17492 1.244
R17824 VSS.n17500 VSS.n17499 1.244
R17825 VSS.n17481 VSS.n17480 1.244
R17826 VSS.n17488 VSS.n17487 1.244
R17827 VSS.n17470 VSS.n17469 1.244
R17828 VSS.n17477 VSS 1.244
R17829 VSS.n17472 VSS.n17471 1.244
R17830 VSS.n17457 VSS.n17456 1.244
R17831 VSS.n17464 VSS.n17463 1.244
R17832 VSS.n17445 VSS.n17444 1.244
R17833 VSS.n17452 VSS.n17451 1.244
R17834 VSS.n17433 VSS.n17432 1.244
R17835 VSS.n17440 VSS.n17439 1.244
R17836 VSS.n17361 VSS.n17360 1.244
R17837 VSS.n17415 VSS.n17414 1.244
R17838 VSS.n17349 VSS.n17348 1.244
R17839 VSS.n17356 VSS.n17355 1.244
R17840 VSS.n17337 VSS.n17336 1.244
R17841 VSS.n17344 VSS.n17343 1.244
R17842 VSS.n17325 VSS.n17324 1.244
R17843 VSS.n17332 VSS.n17331 1.244
R17844 VSS.n17313 VSS.n17312 1.244
R17845 VSS.n17320 VSS.n17319 1.244
R17846 VSS.n17302 VSS.n17301 1.244
R17847 VSS.n17309 VSS 1.244
R17848 VSS.n17304 VSS.n17303 1.244
R17849 VSS.n17289 VSS.n17288 1.244
R17850 VSS.n17296 VSS.n17295 1.244
R17851 VSS.n17277 VSS.n17276 1.244
R17852 VSS.n17284 VSS.n17283 1.244
R17853 VSS.n17265 VSS.n17264 1.244
R17854 VSS.n17272 VSS.n17271 1.244
R17855 VSS.n17193 VSS.n17192 1.244
R17856 VSS.n17247 VSS.n17246 1.244
R17857 VSS.n17181 VSS.n17180 1.244
R17858 VSS.n17188 VSS.n17187 1.244
R17859 VSS.n17169 VSS.n17168 1.244
R17860 VSS.n17176 VSS.n17175 1.244
R17861 VSS.n17157 VSS.n17156 1.244
R17862 VSS.n17164 VSS.n17163 1.244
R17863 VSS.n17145 VSS.n17144 1.244
R17864 VSS.n17152 VSS.n17151 1.244
R17865 VSS.n17134 VSS.n17133 1.244
R17866 VSS.n17141 VSS 1.244
R17867 VSS.n17136 VSS.n17135 1.244
R17868 VSS.n17121 VSS.n17120 1.244
R17869 VSS.n17128 VSS.n17127 1.244
R17870 VSS.n17109 VSS.n17108 1.244
R17871 VSS.n17116 VSS.n17115 1.244
R17872 VSS.n17097 VSS.n17096 1.244
R17873 VSS.n17104 VSS.n17103 1.244
R17874 VSS.n17025 VSS.n17024 1.244
R17875 VSS.n17079 VSS.n17078 1.244
R17876 VSS.n17013 VSS.n17012 1.244
R17877 VSS.n17020 VSS.n17019 1.244
R17878 VSS.n17001 VSS.n17000 1.244
R17879 VSS.n17008 VSS.n17007 1.244
R17880 VSS.n16989 VSS.n16988 1.244
R17881 VSS.n16996 VSS.n16995 1.244
R17882 VSS.n16977 VSS.n16976 1.244
R17883 VSS.n16984 VSS.n16983 1.244
R17884 VSS.n16966 VSS.n16965 1.244
R17885 VSS.n16973 VSS 1.244
R17886 VSS.n16968 VSS.n16967 1.244
R17887 VSS.n16953 VSS.n16952 1.244
R17888 VSS.n16960 VSS.n16959 1.244
R17889 VSS.n16941 VSS.n16940 1.244
R17890 VSS.n16948 VSS.n16947 1.244
R17891 VSS.n16929 VSS.n16928 1.244
R17892 VSS.n16936 VSS.n16935 1.244
R17893 VSS.n16857 VSS.n16856 1.244
R17894 VSS.n16911 VSS.n16910 1.244
R17895 VSS.n16845 VSS.n16844 1.244
R17896 VSS.n16852 VSS.n16851 1.244
R17897 VSS.n16833 VSS.n16832 1.244
R17898 VSS.n16840 VSS.n16839 1.244
R17899 VSS.n16821 VSS.n16820 1.244
R17900 VSS.n16828 VSS.n16827 1.244
R17901 VSS.n16809 VSS.n16808 1.244
R17902 VSS.n16816 VSS.n16815 1.244
R17903 VSS.n16798 VSS.n16797 1.244
R17904 VSS.n16805 VSS 1.244
R17905 VSS.n16800 VSS.n16799 1.244
R17906 VSS.n16785 VSS.n16784 1.244
R17907 VSS.n16792 VSS.n16791 1.244
R17908 VSS.n16773 VSS.n16772 1.244
R17909 VSS.n16780 VSS.n16779 1.244
R17910 VSS.n16761 VSS.n16760 1.244
R17911 VSS.n16768 VSS.n16767 1.244
R17912 VSS.n16689 VSS.n16688 1.244
R17913 VSS.n16743 VSS.n16742 1.244
R17914 VSS.n16677 VSS.n16676 1.244
R17915 VSS.n16684 VSS.n16683 1.244
R17916 VSS.n16665 VSS.n16664 1.244
R17917 VSS.n16672 VSS.n16671 1.244
R17918 VSS.n16653 VSS.n16652 1.244
R17919 VSS.n16660 VSS.n16659 1.244
R17920 VSS.n16641 VSS.n16640 1.244
R17921 VSS.n16648 VSS.n16647 1.244
R17922 VSS.n16630 VSS.n16629 1.244
R17923 VSS.n16637 VSS 1.244
R17924 VSS.n16632 VSS.n16631 1.244
R17925 VSS.n16617 VSS.n16616 1.244
R17926 VSS.n16624 VSS.n16623 1.244
R17927 VSS.n16605 VSS.n16604 1.244
R17928 VSS.n16612 VSS.n16611 1.244
R17929 VSS.n16593 VSS.n16592 1.244
R17930 VSS.n16600 VSS.n16599 1.244
R17931 VSS.n13912 VSS.n13911 1.244
R17932 VSS.n13919 VSS.n13918 1.244
R17933 VSS.n13924 VSS.n13923 1.244
R17934 VSS.n13931 VSS.n13930 1.244
R17935 VSS.n13936 VSS.n13935 1.244
R17936 VSS.n13943 VSS.n13942 1.244
R17937 VSS.n13948 VSS.n13947 1.244
R17938 VSS.n13955 VSS.n13954 1.244
R17939 VSS.n13960 VSS.n13959 1.244
R17940 VSS.n13967 VSS.n13966 1.244
R17941 VSS.n13972 VSS.n13971 1.244
R17942 VSS VSS.n13977 1.244
R17943 VSS.n13979 VSS.n13978 1.244
R17944 VSS.n13984 VSS.n13983 1.244
R17945 VSS.n13991 VSS.n13990 1.244
R17946 VSS.n13996 VSS.n13995 1.244
R17947 VSS.n14003 VSS.n14002 1.244
R17948 VSS.n14008 VSS.n14007 1.244
R17949 VSS.n14060 VSS.n14059 1.244
R17950 VSS.n13732 VSS.n13731 1.244
R17951 VSS.n13739 VSS.n13738 1.244
R17952 VSS.n13744 VSS.n13743 1.244
R17953 VSS.n13751 VSS.n13750 1.244
R17954 VSS.n13756 VSS.n13755 1.244
R17955 VSS.n13763 VSS.n13762 1.244
R17956 VSS.n13768 VSS.n13767 1.244
R17957 VSS.n13775 VSS.n13774 1.244
R17958 VSS.n13780 VSS.n13779 1.244
R17959 VSS.n13787 VSS.n13786 1.244
R17960 VSS.n13792 VSS.n13791 1.244
R17961 VSS VSS.n13797 1.244
R17962 VSS.n13799 VSS.n13798 1.244
R17963 VSS.n13804 VSS.n13803 1.244
R17964 VSS.n13811 VSS.n13810 1.244
R17965 VSS.n13816 VSS.n13815 1.244
R17966 VSS.n13823 VSS.n13822 1.244
R17967 VSS.n13828 VSS.n13827 1.244
R17968 VSS.n13880 VSS.n13879 1.244
R17969 VSS.n13552 VSS.n13551 1.244
R17970 VSS.n13559 VSS.n13558 1.244
R17971 VSS.n13564 VSS.n13563 1.244
R17972 VSS.n13571 VSS.n13570 1.244
R17973 VSS.n13576 VSS.n13575 1.244
R17974 VSS.n13583 VSS.n13582 1.244
R17975 VSS.n13588 VSS.n13587 1.244
R17976 VSS.n13595 VSS.n13594 1.244
R17977 VSS.n13600 VSS.n13599 1.244
R17978 VSS.n13607 VSS.n13606 1.244
R17979 VSS.n13612 VSS.n13611 1.244
R17980 VSS VSS.n13617 1.244
R17981 VSS.n13619 VSS.n13618 1.244
R17982 VSS.n13624 VSS.n13623 1.244
R17983 VSS.n13631 VSS.n13630 1.244
R17984 VSS.n13636 VSS.n13635 1.244
R17985 VSS.n13643 VSS.n13642 1.244
R17986 VSS.n13648 VSS.n13647 1.244
R17987 VSS.n13700 VSS.n13699 1.244
R17988 VSS.n13372 VSS.n13371 1.244
R17989 VSS.n13379 VSS.n13378 1.244
R17990 VSS.n13384 VSS.n13383 1.244
R17991 VSS.n13391 VSS.n13390 1.244
R17992 VSS.n13396 VSS.n13395 1.244
R17993 VSS.n13403 VSS.n13402 1.244
R17994 VSS.n13408 VSS.n13407 1.244
R17995 VSS.n13415 VSS.n13414 1.244
R17996 VSS.n13420 VSS.n13419 1.244
R17997 VSS.n13427 VSS.n13426 1.244
R17998 VSS.n13432 VSS.n13431 1.244
R17999 VSS VSS.n13437 1.244
R18000 VSS.n13439 VSS.n13438 1.244
R18001 VSS.n13444 VSS.n13443 1.244
R18002 VSS.n13451 VSS.n13450 1.244
R18003 VSS.n13456 VSS.n13455 1.244
R18004 VSS.n13463 VSS.n13462 1.244
R18005 VSS.n13468 VSS.n13467 1.244
R18006 VSS.n13520 VSS.n13519 1.244
R18007 VSS.n13192 VSS.n13191 1.244
R18008 VSS.n13199 VSS.n13198 1.244
R18009 VSS.n13204 VSS.n13203 1.244
R18010 VSS.n13211 VSS.n13210 1.244
R18011 VSS.n13216 VSS.n13215 1.244
R18012 VSS.n13223 VSS.n13222 1.244
R18013 VSS.n13228 VSS.n13227 1.244
R18014 VSS.n13235 VSS.n13234 1.244
R18015 VSS.n13240 VSS.n13239 1.244
R18016 VSS.n13247 VSS.n13246 1.244
R18017 VSS.n13252 VSS.n13251 1.244
R18018 VSS VSS.n13257 1.244
R18019 VSS.n13259 VSS.n13258 1.244
R18020 VSS.n13264 VSS.n13263 1.244
R18021 VSS.n13271 VSS.n13270 1.244
R18022 VSS.n13276 VSS.n13275 1.244
R18023 VSS.n13283 VSS.n13282 1.244
R18024 VSS.n13288 VSS.n13287 1.244
R18025 VSS.n13340 VSS.n13339 1.244
R18026 VSS.n13012 VSS.n13011 1.244
R18027 VSS.n13019 VSS.n13018 1.244
R18028 VSS.n13024 VSS.n13023 1.244
R18029 VSS.n13031 VSS.n13030 1.244
R18030 VSS.n13036 VSS.n13035 1.244
R18031 VSS.n13043 VSS.n13042 1.244
R18032 VSS.n13048 VSS.n13047 1.244
R18033 VSS.n13055 VSS.n13054 1.244
R18034 VSS.n13060 VSS.n13059 1.244
R18035 VSS.n13067 VSS.n13066 1.244
R18036 VSS.n13072 VSS.n13071 1.244
R18037 VSS VSS.n13077 1.244
R18038 VSS.n13079 VSS.n13078 1.244
R18039 VSS.n13084 VSS.n13083 1.244
R18040 VSS.n13091 VSS.n13090 1.244
R18041 VSS.n13096 VSS.n13095 1.244
R18042 VSS.n13103 VSS.n13102 1.244
R18043 VSS.n13108 VSS.n13107 1.244
R18044 VSS.n13160 VSS.n13159 1.244
R18045 VSS.n12832 VSS.n12831 1.244
R18046 VSS.n12839 VSS.n12838 1.244
R18047 VSS.n12844 VSS.n12843 1.244
R18048 VSS.n12851 VSS.n12850 1.244
R18049 VSS.n12856 VSS.n12855 1.244
R18050 VSS.n12863 VSS.n12862 1.244
R18051 VSS.n12868 VSS.n12867 1.244
R18052 VSS.n12875 VSS.n12874 1.244
R18053 VSS.n12880 VSS.n12879 1.244
R18054 VSS.n12887 VSS.n12886 1.244
R18055 VSS.n12892 VSS.n12891 1.244
R18056 VSS VSS.n12897 1.244
R18057 VSS.n12899 VSS.n12898 1.244
R18058 VSS.n12904 VSS.n12903 1.244
R18059 VSS.n12911 VSS.n12910 1.244
R18060 VSS.n12916 VSS.n12915 1.244
R18061 VSS.n12923 VSS.n12922 1.244
R18062 VSS.n12928 VSS.n12927 1.244
R18063 VSS.n12980 VSS.n12979 1.244
R18064 VSS.n12652 VSS.n12651 1.244
R18065 VSS.n12659 VSS.n12658 1.244
R18066 VSS.n12664 VSS.n12663 1.244
R18067 VSS.n12671 VSS.n12670 1.244
R18068 VSS.n12676 VSS.n12675 1.244
R18069 VSS.n12683 VSS.n12682 1.244
R18070 VSS.n12688 VSS.n12687 1.244
R18071 VSS.n12695 VSS.n12694 1.244
R18072 VSS.n12700 VSS.n12699 1.244
R18073 VSS.n12707 VSS.n12706 1.244
R18074 VSS.n12712 VSS.n12711 1.244
R18075 VSS VSS.n12717 1.244
R18076 VSS.n12719 VSS.n12718 1.244
R18077 VSS.n12724 VSS.n12723 1.244
R18078 VSS.n12731 VSS.n12730 1.244
R18079 VSS.n12736 VSS.n12735 1.244
R18080 VSS.n12743 VSS.n12742 1.244
R18081 VSS.n12748 VSS.n12747 1.244
R18082 VSS.n12800 VSS.n12799 1.244
R18083 VSS.n9319 VSS.n9318 1.244
R18084 VSS.n9371 VSS.n9370 1.244
R18085 VSS.n9307 VSS.n9306 1.244
R18086 VSS.n9314 VSS.n9313 1.244
R18087 VSS.n9295 VSS.n9294 1.244
R18088 VSS.n9302 VSS.n9301 1.244
R18089 VSS.n9283 VSS.n9282 1.244
R18090 VSS.n9290 VSS.n9289 1.244
R18091 VSS.n9271 VSS.n9270 1.244
R18092 VSS.n9278 VSS.n9277 1.244
R18093 VSS.n9260 VSS.n9259 1.244
R18094 VSS.n9267 VSS 1.244
R18095 VSS.n9262 VSS.n9261 1.244
R18096 VSS.n9247 VSS.n9246 1.244
R18097 VSS.n9254 VSS.n9253 1.244
R18098 VSS.n9235 VSS.n9234 1.244
R18099 VSS.n9242 VSS.n9241 1.244
R18100 VSS.n9223 VSS.n9222 1.244
R18101 VSS.n9230 VSS.n9229 1.244
R18102 VSS.n9487 VSS.n9486 1.244
R18103 VSS.n9539 VSS.n9538 1.244
R18104 VSS.n9475 VSS.n9474 1.244
R18105 VSS.n9482 VSS.n9481 1.244
R18106 VSS.n9463 VSS.n9462 1.244
R18107 VSS.n9470 VSS.n9469 1.244
R18108 VSS.n9451 VSS.n9450 1.244
R18109 VSS.n9458 VSS.n9457 1.244
R18110 VSS.n9439 VSS.n9438 1.244
R18111 VSS.n9446 VSS.n9445 1.244
R18112 VSS.n9428 VSS.n9427 1.244
R18113 VSS.n9435 VSS 1.244
R18114 VSS.n9430 VSS.n9429 1.244
R18115 VSS.n9415 VSS.n9414 1.244
R18116 VSS.n9422 VSS.n9421 1.244
R18117 VSS.n9403 VSS.n9402 1.244
R18118 VSS.n9410 VSS.n9409 1.244
R18119 VSS.n9391 VSS.n9390 1.244
R18120 VSS.n9398 VSS.n9397 1.244
R18121 VSS.n9655 VSS.n9654 1.244
R18122 VSS.n9707 VSS.n9706 1.244
R18123 VSS.n9643 VSS.n9642 1.244
R18124 VSS.n9650 VSS.n9649 1.244
R18125 VSS.n9631 VSS.n9630 1.244
R18126 VSS.n9638 VSS.n9637 1.244
R18127 VSS.n9619 VSS.n9618 1.244
R18128 VSS.n9626 VSS.n9625 1.244
R18129 VSS.n9607 VSS.n9606 1.244
R18130 VSS.n9614 VSS.n9613 1.244
R18131 VSS.n9596 VSS.n9595 1.244
R18132 VSS.n9603 VSS 1.244
R18133 VSS.n9598 VSS.n9597 1.244
R18134 VSS.n9583 VSS.n9582 1.244
R18135 VSS.n9590 VSS.n9589 1.244
R18136 VSS.n9571 VSS.n9570 1.244
R18137 VSS.n9578 VSS.n9577 1.244
R18138 VSS.n9559 VSS.n9558 1.244
R18139 VSS.n9566 VSS.n9565 1.244
R18140 VSS.n9823 VSS.n9822 1.244
R18141 VSS.n9875 VSS.n9874 1.244
R18142 VSS.n9811 VSS.n9810 1.244
R18143 VSS.n9818 VSS.n9817 1.244
R18144 VSS.n9799 VSS.n9798 1.244
R18145 VSS.n9806 VSS.n9805 1.244
R18146 VSS.n9787 VSS.n9786 1.244
R18147 VSS.n9794 VSS.n9793 1.244
R18148 VSS.n9775 VSS.n9774 1.244
R18149 VSS.n9782 VSS.n9781 1.244
R18150 VSS.n9764 VSS.n9763 1.244
R18151 VSS.n9771 VSS 1.244
R18152 VSS.n9766 VSS.n9765 1.244
R18153 VSS.n9751 VSS.n9750 1.244
R18154 VSS.n9758 VSS.n9757 1.244
R18155 VSS.n9739 VSS.n9738 1.244
R18156 VSS.n9746 VSS.n9745 1.244
R18157 VSS.n9727 VSS.n9726 1.244
R18158 VSS.n9734 VSS.n9733 1.244
R18159 VSS.n9991 VSS.n9990 1.244
R18160 VSS.n10043 VSS.n10042 1.244
R18161 VSS.n9979 VSS.n9978 1.244
R18162 VSS.n9986 VSS.n9985 1.244
R18163 VSS.n9967 VSS.n9966 1.244
R18164 VSS.n9974 VSS.n9973 1.244
R18165 VSS.n9955 VSS.n9954 1.244
R18166 VSS.n9962 VSS.n9961 1.244
R18167 VSS.n9943 VSS.n9942 1.244
R18168 VSS.n9950 VSS.n9949 1.244
R18169 VSS.n9932 VSS.n9931 1.244
R18170 VSS.n9939 VSS 1.244
R18171 VSS.n9934 VSS.n9933 1.244
R18172 VSS.n9919 VSS.n9918 1.244
R18173 VSS.n9926 VSS.n9925 1.244
R18174 VSS.n9907 VSS.n9906 1.244
R18175 VSS.n9914 VSS.n9913 1.244
R18176 VSS.n9895 VSS.n9894 1.244
R18177 VSS.n9902 VSS.n9901 1.244
R18178 VSS.n10159 VSS.n10158 1.244
R18179 VSS.n10211 VSS.n10210 1.244
R18180 VSS.n10147 VSS.n10146 1.244
R18181 VSS.n10154 VSS.n10153 1.244
R18182 VSS.n10135 VSS.n10134 1.244
R18183 VSS.n10142 VSS.n10141 1.244
R18184 VSS.n10123 VSS.n10122 1.244
R18185 VSS.n10130 VSS.n10129 1.244
R18186 VSS.n10111 VSS.n10110 1.244
R18187 VSS.n10118 VSS.n10117 1.244
R18188 VSS.n10100 VSS.n10099 1.244
R18189 VSS.n10107 VSS 1.244
R18190 VSS.n10102 VSS.n10101 1.244
R18191 VSS.n10087 VSS.n10086 1.244
R18192 VSS.n10094 VSS.n10093 1.244
R18193 VSS.n10075 VSS.n10074 1.244
R18194 VSS.n10082 VSS.n10081 1.244
R18195 VSS.n10063 VSS.n10062 1.244
R18196 VSS.n10070 VSS.n10069 1.244
R18197 VSS.n10327 VSS.n10326 1.244
R18198 VSS.n10379 VSS.n10378 1.244
R18199 VSS.n10315 VSS.n10314 1.244
R18200 VSS.n10322 VSS.n10321 1.244
R18201 VSS.n10303 VSS.n10302 1.244
R18202 VSS.n10310 VSS.n10309 1.244
R18203 VSS.n10291 VSS.n10290 1.244
R18204 VSS.n10298 VSS.n10297 1.244
R18205 VSS.n10279 VSS.n10278 1.244
R18206 VSS.n10286 VSS.n10285 1.244
R18207 VSS.n10268 VSS.n10267 1.244
R18208 VSS.n10275 VSS 1.244
R18209 VSS.n10270 VSS.n10269 1.244
R18210 VSS.n10255 VSS.n10254 1.244
R18211 VSS.n10262 VSS.n10261 1.244
R18212 VSS.n10243 VSS.n10242 1.244
R18213 VSS.n10250 VSS.n10249 1.244
R18214 VSS.n10231 VSS.n10230 1.244
R18215 VSS.n10238 VSS.n10237 1.244
R18216 VSS.n10494 VSS.n10493 1.244
R18217 VSS.n10547 VSS.n10546 1.244
R18218 VSS.n10482 VSS.n10481 1.244
R18219 VSS.n10489 VSS.n10488 1.244
R18220 VSS.n10470 VSS.n10469 1.244
R18221 VSS.n10477 VSS.n10476 1.244
R18222 VSS.n10458 VSS.n10457 1.244
R18223 VSS.n10465 VSS.n10464 1.244
R18224 VSS.n10446 VSS.n10445 1.244
R18225 VSS.n10453 VSS.n10452 1.244
R18226 VSS.n10435 VSS.n10434 1.244
R18227 VSS.n10442 VSS 1.244
R18228 VSS.n10437 VSS.n10436 1.244
R18229 VSS.n10422 VSS.n10421 1.244
R18230 VSS.n10429 VSS.n10428 1.244
R18231 VSS.n10410 VSS.n10409 1.244
R18232 VSS.n10417 VSS.n10416 1.244
R18233 VSS.n10398 VSS.n10397 1.244
R18234 VSS.n10405 VSS.n10404 1.244
R18235 VSS.n2378 VSS.n2377 1.244
R18236 VSS.n2380 VSS.n2324 1.244
R18237 VSS.n2455 VSS.n2454 1.244
R18238 VSS.n2448 VSS.n2325 1.244
R18239 VSS.n2447 VSS.n2445 1.244
R18240 VSS.n2442 VSS.n2384 1.244
R18241 VSS.n2388 VSS.n2387 1.244
R18242 VSS.n2436 VSS.n2435 1.244
R18243 VSS.n2392 VSS.n2390 1.244
R18244 VSS.n2430 VSS.n2429 1.244
R18245 VSS.n2396 VSS.n2394 1.244
R18246 VSS.n2426 VSS 1.244
R18247 VSS.n2424 VSS.n2423 1.244
R18248 VSS.n2397 VSS.n2314 1.244
R18249 VSS.n2419 VSS.n2418 1.244
R18250 VSS.n2402 VSS.n2400 1.244
R18251 VSS.n2413 VSS.n2412 1.244
R18252 VSS.n2407 VSS.n2403 1.244
R18253 VSS.n2408 VSS.n2286 1.244
R18254 VSS.n2468 VSS.n2467 1.244
R18255 VSS.n2470 VSS.n2234 1.244
R18256 VSS.n2545 VSS.n2544 1.244
R18257 VSS.n2538 VSS.n2235 1.244
R18258 VSS.n2537 VSS.n2535 1.244
R18259 VSS.n2532 VSS.n2474 1.244
R18260 VSS.n2478 VSS.n2477 1.244
R18261 VSS.n2526 VSS.n2525 1.244
R18262 VSS.n2482 VSS.n2480 1.244
R18263 VSS.n2520 VSS.n2519 1.244
R18264 VSS.n2486 VSS.n2484 1.244
R18265 VSS.n2516 VSS 1.244
R18266 VSS.n2514 VSS.n2513 1.244
R18267 VSS.n2487 VSS.n2224 1.244
R18268 VSS.n2509 VSS.n2508 1.244
R18269 VSS.n2492 VSS.n2490 1.244
R18270 VSS.n2503 VSS.n2502 1.244
R18271 VSS.n2497 VSS.n2493 1.244
R18272 VSS.n2498 VSS.n2196 1.244
R18273 VSS.n2558 VSS.n2557 1.244
R18274 VSS.n2560 VSS.n2144 1.244
R18275 VSS.n2635 VSS.n2634 1.244
R18276 VSS.n2628 VSS.n2145 1.244
R18277 VSS.n2627 VSS.n2625 1.244
R18278 VSS.n2622 VSS.n2564 1.244
R18279 VSS.n2568 VSS.n2567 1.244
R18280 VSS.n2616 VSS.n2615 1.244
R18281 VSS.n2572 VSS.n2570 1.244
R18282 VSS.n2610 VSS.n2609 1.244
R18283 VSS.n2576 VSS.n2574 1.244
R18284 VSS.n2606 VSS 1.244
R18285 VSS.n2604 VSS.n2603 1.244
R18286 VSS.n2577 VSS.n2134 1.244
R18287 VSS.n2599 VSS.n2598 1.244
R18288 VSS.n2582 VSS.n2580 1.244
R18289 VSS.n2593 VSS.n2592 1.244
R18290 VSS.n2587 VSS.n2583 1.244
R18291 VSS.n2588 VSS.n2106 1.244
R18292 VSS.n2648 VSS.n2647 1.244
R18293 VSS.n2650 VSS.n2054 1.244
R18294 VSS.n2725 VSS.n2724 1.244
R18295 VSS.n2718 VSS.n2055 1.244
R18296 VSS.n2717 VSS.n2715 1.244
R18297 VSS.n2712 VSS.n2654 1.244
R18298 VSS.n2658 VSS.n2657 1.244
R18299 VSS.n2706 VSS.n2705 1.244
R18300 VSS.n2662 VSS.n2660 1.244
R18301 VSS.n2700 VSS.n2699 1.244
R18302 VSS.n2666 VSS.n2664 1.244
R18303 VSS.n2696 VSS 1.244
R18304 VSS.n2694 VSS.n2693 1.244
R18305 VSS.n2667 VSS.n2044 1.244
R18306 VSS.n2689 VSS.n2688 1.244
R18307 VSS.n2672 VSS.n2670 1.244
R18308 VSS.n2683 VSS.n2682 1.244
R18309 VSS.n2677 VSS.n2673 1.244
R18310 VSS.n2678 VSS.n2016 1.244
R18311 VSS.n2738 VSS.n2737 1.244
R18312 VSS.n2740 VSS.n1964 1.244
R18313 VSS.n2815 VSS.n2814 1.244
R18314 VSS.n2808 VSS.n1965 1.244
R18315 VSS.n2807 VSS.n2805 1.244
R18316 VSS.n2802 VSS.n2744 1.244
R18317 VSS.n2748 VSS.n2747 1.244
R18318 VSS.n2796 VSS.n2795 1.244
R18319 VSS.n2752 VSS.n2750 1.244
R18320 VSS.n2790 VSS.n2789 1.244
R18321 VSS.n2756 VSS.n2754 1.244
R18322 VSS.n2786 VSS 1.244
R18323 VSS.n2784 VSS.n2783 1.244
R18324 VSS.n2757 VSS.n1954 1.244
R18325 VSS.n2779 VSS.n2778 1.244
R18326 VSS.n2762 VSS.n2760 1.244
R18327 VSS.n2773 VSS.n2772 1.244
R18328 VSS.n2767 VSS.n2763 1.244
R18329 VSS.n2768 VSS.n1926 1.244
R18330 VSS.n2828 VSS.n2827 1.244
R18331 VSS.n2830 VSS.n1874 1.244
R18332 VSS.n2905 VSS.n2904 1.244
R18333 VSS.n2898 VSS.n1875 1.244
R18334 VSS.n2897 VSS.n2895 1.244
R18335 VSS.n2892 VSS.n2834 1.244
R18336 VSS.n2838 VSS.n2837 1.244
R18337 VSS.n2886 VSS.n2885 1.244
R18338 VSS.n2842 VSS.n2840 1.244
R18339 VSS.n2880 VSS.n2879 1.244
R18340 VSS.n2846 VSS.n2844 1.244
R18341 VSS.n2876 VSS 1.244
R18342 VSS.n2874 VSS.n2873 1.244
R18343 VSS.n2847 VSS.n1864 1.244
R18344 VSS.n2869 VSS.n2868 1.244
R18345 VSS.n2852 VSS.n2850 1.244
R18346 VSS.n2863 VSS.n2862 1.244
R18347 VSS.n2857 VSS.n2853 1.244
R18348 VSS.n2858 VSS.n1836 1.244
R18349 VSS.n2918 VSS.n2917 1.244
R18350 VSS.n2920 VSS.n1784 1.244
R18351 VSS.n2995 VSS.n2994 1.244
R18352 VSS.n2988 VSS.n1785 1.244
R18353 VSS.n2987 VSS.n2985 1.244
R18354 VSS.n2982 VSS.n2924 1.244
R18355 VSS.n2928 VSS.n2927 1.244
R18356 VSS.n2976 VSS.n2975 1.244
R18357 VSS.n2932 VSS.n2930 1.244
R18358 VSS.n2970 VSS.n2969 1.244
R18359 VSS.n2936 VSS.n2934 1.244
R18360 VSS.n2966 VSS 1.244
R18361 VSS.n2964 VSS.n2963 1.244
R18362 VSS.n2937 VSS.n1774 1.244
R18363 VSS.n2959 VSS.n2958 1.244
R18364 VSS.n2942 VSS.n2940 1.244
R18365 VSS.n2953 VSS.n2952 1.244
R18366 VSS.n2947 VSS.n2943 1.244
R18367 VSS.n2948 VSS.n1746 1.244
R18368 VSS.n3008 VSS.n3007 1.244
R18369 VSS.n3010 VSS.n1694 1.244
R18370 VSS.n3085 VSS.n3084 1.244
R18371 VSS.n3078 VSS.n1695 1.244
R18372 VSS.n3077 VSS.n3075 1.244
R18373 VSS.n3072 VSS.n3014 1.244
R18374 VSS.n3018 VSS.n3017 1.244
R18375 VSS.n3066 VSS.n3065 1.244
R18376 VSS.n3022 VSS.n3020 1.244
R18377 VSS.n3060 VSS.n3059 1.244
R18378 VSS.n3026 VSS.n3024 1.244
R18379 VSS.n3056 VSS 1.244
R18380 VSS.n3054 VSS.n3053 1.244
R18381 VSS.n3027 VSS.n1684 1.244
R18382 VSS.n3049 VSS.n3048 1.244
R18383 VSS.n3032 VSS.n3030 1.244
R18384 VSS.n3043 VSS.n3042 1.244
R18385 VSS.n3037 VSS.n3033 1.244
R18386 VSS.n3038 VSS.n1656 1.244
R18387 VSS.n6250 VSS.n6075 1.244
R18388 VSS.n6131 VSS.n6128 1.244
R18389 VSS.n6130 VSS.n6124 1.244
R18390 VSS.n6139 VSS.n6136 1.244
R18391 VSS.n6138 VSS.n6122 1.244
R18392 VSS.n6147 VSS.n6144 1.244
R18393 VSS.n6146 VSS.n6120 1.244
R18394 VSS.n6155 VSS.n6152 1.244
R18395 VSS.n6154 VSS.n6118 1.244
R18396 VSS.n6163 VSS.n6160 1.244
R18397 VSS.n6162 VSS.n6116 1.244
R18398 VSS VSS.n6167 1.244
R18399 VSS.n6171 VSS.n6168 1.244
R18400 VSS.n6170 VSS.n6114 1.244
R18401 VSS.n6179 VSS.n6176 1.244
R18402 VSS.n6178 VSS.n6112 1.244
R18403 VSS.n6187 VSS.n6184 1.244
R18404 VSS.n6186 VSS.n6109 1.244
R18405 VSS.n6241 VSS.n6110 1.244
R18406 VSS.n6314 VSS.n5959 1.244
R18407 VSS.n6015 VSS.n6012 1.244
R18408 VSS.n6014 VSS.n6008 1.244
R18409 VSS.n6023 VSS.n6020 1.244
R18410 VSS.n6022 VSS.n6006 1.244
R18411 VSS.n6031 VSS.n6028 1.244
R18412 VSS.n6030 VSS.n6004 1.244
R18413 VSS.n6039 VSS.n6036 1.244
R18414 VSS.n6038 VSS.n6002 1.244
R18415 VSS.n6047 VSS.n6044 1.244
R18416 VSS.n6046 VSS.n6000 1.244
R18417 VSS VSS.n6051 1.244
R18418 VSS.n6055 VSS.n6052 1.244
R18419 VSS.n6054 VSS.n5998 1.244
R18420 VSS.n6063 VSS.n6060 1.244
R18421 VSS.n6062 VSS.n5996 1.244
R18422 VSS.n6071 VSS.n6068 1.244
R18423 VSS.n6070 VSS.n5993 1.244
R18424 VSS.n6305 VSS.n5994 1.244
R18425 VSS.n6378 VSS.n5843 1.244
R18426 VSS.n5899 VSS.n5896 1.244
R18427 VSS.n5898 VSS.n5892 1.244
R18428 VSS.n5907 VSS.n5904 1.244
R18429 VSS.n5906 VSS.n5890 1.244
R18430 VSS.n5915 VSS.n5912 1.244
R18431 VSS.n5914 VSS.n5888 1.244
R18432 VSS.n5923 VSS.n5920 1.244
R18433 VSS.n5922 VSS.n5886 1.244
R18434 VSS.n5931 VSS.n5928 1.244
R18435 VSS.n5930 VSS.n5884 1.244
R18436 VSS VSS.n5935 1.244
R18437 VSS.n5939 VSS.n5936 1.244
R18438 VSS.n5938 VSS.n5882 1.244
R18439 VSS.n5947 VSS.n5944 1.244
R18440 VSS.n5946 VSS.n5880 1.244
R18441 VSS.n5955 VSS.n5952 1.244
R18442 VSS.n5954 VSS.n5877 1.244
R18443 VSS.n6369 VSS.n5878 1.244
R18444 VSS.n6940 VSS.n5787 1.244
R18445 VSS.n5791 VSS.n5788 1.244
R18446 VSS.n7039 VSS.n7038 1.244
R18447 VSS.n5796 VSS.n5792 1.244
R18448 VSS.n7033 VSS.n7032 1.244
R18449 VSS.n5802 VSS.n5797 1.244
R18450 VSS.n7027 VSS.n7026 1.244
R18451 VSS.n5808 VSS.n5803 1.244
R18452 VSS.n7021 VSS.n7020 1.244
R18453 VSS.n5814 VSS.n5809 1.244
R18454 VSS.n7015 VSS.n7014 1.244
R18455 VSS.n7013 VSS 1.244
R18456 VSS.n5821 VSS.n5819 1.244
R18457 VSS.n7009 VSS.n7008 1.244
R18458 VSS.n5826 VSS.n5820 1.244
R18459 VSS.n7003 VSS.n7002 1.244
R18460 VSS.n5832 VSS.n5827 1.244
R18461 VSS.n6997 VSS.n6996 1.244
R18462 VSS.n5838 VSS.n5833 1.244
R18463 VSS.n6852 VSS.n6850 1.244
R18464 VSS.n6854 VSS.n6438 1.244
R18465 VSS.n6928 VSS.n6927 1.244
R18466 VSS.n6921 VSS.n6439 1.244
R18467 VSS.n6920 VSS.n6918 1.244
R18468 VSS.n6915 VSS.n6858 1.244
R18469 VSS.n6862 VSS.n6861 1.244
R18470 VSS.n6909 VSS.n6908 1.244
R18471 VSS.n6866 VSS.n6864 1.244
R18472 VSS.n6903 VSS.n6902 1.244
R18473 VSS.n6870 VSS.n6868 1.244
R18474 VSS.n6899 VSS 1.244
R18475 VSS.n6897 VSS.n6896 1.244
R18476 VSS.n6874 VSS.n6872 1.244
R18477 VSS.n6891 VSS.n6890 1.244
R18478 VSS.n6875 VSS.n6428 1.244
R18479 VSS.n6886 VSS.n6885 1.244
R18480 VSS.n6880 VSS.n6878 1.244
R18481 VSS.n6881 VSS.n6400 1.244
R18482 VSS.n6762 VSS.n6760 1.244
R18483 VSS.n6764 VSS.n6528 1.244
R18484 VSS.n6838 VSS.n6837 1.244
R18485 VSS.n6831 VSS.n6529 1.244
R18486 VSS.n6830 VSS.n6828 1.244
R18487 VSS.n6825 VSS.n6768 1.244
R18488 VSS.n6772 VSS.n6771 1.244
R18489 VSS.n6819 VSS.n6818 1.244
R18490 VSS.n6776 VSS.n6774 1.244
R18491 VSS.n6813 VSS.n6812 1.244
R18492 VSS.n6780 VSS.n6778 1.244
R18493 VSS.n6809 VSS 1.244
R18494 VSS.n6807 VSS.n6806 1.244
R18495 VSS.n6784 VSS.n6782 1.244
R18496 VSS.n6801 VSS.n6800 1.244
R18497 VSS.n6785 VSS.n6518 1.244
R18498 VSS.n6796 VSS.n6795 1.244
R18499 VSS.n6790 VSS.n6788 1.244
R18500 VSS.n6791 VSS.n6490 1.244
R18501 VSS.n6672 VSS.n6670 1.244
R18502 VSS.n6674 VSS.n6618 1.244
R18503 VSS.n6748 VSS.n6747 1.244
R18504 VSS.n6741 VSS.n6619 1.244
R18505 VSS.n6740 VSS.n6738 1.244
R18506 VSS.n6735 VSS.n6678 1.244
R18507 VSS.n6682 VSS.n6681 1.244
R18508 VSS.n6729 VSS.n6728 1.244
R18509 VSS.n6686 VSS.n6684 1.244
R18510 VSS.n6723 VSS.n6722 1.244
R18511 VSS.n6690 VSS.n6688 1.244
R18512 VSS.n6719 VSS 1.244
R18513 VSS.n6717 VSS.n6716 1.244
R18514 VSS.n6694 VSS.n6692 1.244
R18515 VSS.n6711 VSS.n6710 1.244
R18516 VSS.n6695 VSS.n6608 1.244
R18517 VSS.n6706 VSS.n6705 1.244
R18518 VSS.n6700 VSS.n6698 1.244
R18519 VSS.n6701 VSS.n6580 1.244
R18520 VSS.n18024 VSS.n18023 1.206
R18521 VSS.n17767 VSS.n17743 1.142
R18522 VSS VSS.n18024 1.07
R18523 VSS.n18020 VSS.n18019 1.065
R18524 VSS.n5133 VSS.n5132 1.01
R18525 VSS.n18024 VSS 0.969
R18526 VSS.n16381 VSS.n16380 0.905
R18527 VSS.n16390 VSS.n16389 0.905
R18528 VSS.n16395 VSS.n16394 0.905
R18529 VSS.n16404 VSS.n16403 0.905
R18530 VSS.n16409 VSS.n16408 0.905
R18531 VSS.n16418 VSS.n16417 0.905
R18532 VSS.n16423 VSS.n16422 0.905
R18533 VSS.n16432 VSS.n16431 0.905
R18534 VSS.n16437 VSS.n16436 0.905
R18535 VSS.n16446 VSS.n16445 0.905
R18536 VSS.n16451 VSS.n16450 0.905
R18537 VSS.n16465 VSS.n16464 0.905
R18538 VSS.n16463 VSS.n14555 0.905
R18539 VSS.n14557 VSS.n14556 0.905
R18540 VSS.n14554 VSS.n14553 0.905
R18541 VSS.n16482 VSS.n16481 0.905
R18542 VSS.n16487 VSS.n16486 0.905
R18543 VSS.n16496 VSS.n16495 0.905
R18544 VSS.n16501 VSS.n16500 0.905
R18545 VSS.n16510 VSS.n16509 0.905
R18546 VSS.n16515 VSS.n16514 0.905
R18547 VSS.n16524 VSS.n16523 0.905
R18548 VSS.n16574 VSS.n16573 0.905
R18549 VSS.n16585 VSS.n16584 0.905
R18550 VSS.n16125 VSS.n16124 0.905
R18551 VSS.n16134 VSS.n16133 0.905
R18552 VSS.n16139 VSS.n16138 0.905
R18553 VSS.n16148 VSS.n16147 0.905
R18554 VSS.n16153 VSS.n16152 0.905
R18555 VSS.n16162 VSS.n16161 0.905
R18556 VSS.n16167 VSS.n16166 0.905
R18557 VSS.n16176 VSS.n16175 0.905
R18558 VSS.n16181 VSS.n16180 0.905
R18559 VSS.n16190 VSS.n16189 0.905
R18560 VSS.n16195 VSS.n16194 0.905
R18561 VSS.n16209 VSS.n16208 0.905
R18562 VSS.n16207 VSS.n14561 0.905
R18563 VSS.n14563 VSS.n14562 0.905
R18564 VSS.n14560 VSS.n14559 0.905
R18565 VSS.n16226 VSS.n16225 0.905
R18566 VSS.n16231 VSS.n16230 0.905
R18567 VSS.n16240 VSS.n16239 0.905
R18568 VSS.n16245 VSS.n16244 0.905
R18569 VSS.n16254 VSS.n16253 0.905
R18570 VSS.n16259 VSS.n16258 0.905
R18571 VSS.n16268 VSS.n16267 0.905
R18572 VSS.n16273 VSS.n16272 0.905
R18573 VSS.n15881 VSS.n15880 0.905
R18574 VSS.n15890 VSS.n15889 0.905
R18575 VSS.n15895 VSS.n15894 0.905
R18576 VSS.n15904 VSS.n15903 0.905
R18577 VSS.n15909 VSS.n15908 0.905
R18578 VSS.n15918 VSS.n15917 0.905
R18579 VSS.n15923 VSS.n15922 0.905
R18580 VSS.n15932 VSS.n15931 0.905
R18581 VSS.n15937 VSS.n15936 0.905
R18582 VSS.n15946 VSS.n15945 0.905
R18583 VSS.n15951 VSS.n15950 0.905
R18584 VSS.n15965 VSS.n15964 0.905
R18585 VSS.n15963 VSS.n14567 0.905
R18586 VSS.n14569 VSS.n14568 0.905
R18587 VSS.n14566 VSS.n14565 0.905
R18588 VSS.n15982 VSS.n15981 0.905
R18589 VSS.n15987 VSS.n15986 0.905
R18590 VSS.n15996 VSS.n15995 0.905
R18591 VSS.n16001 VSS.n16000 0.905
R18592 VSS.n16010 VSS.n16009 0.905
R18593 VSS.n16015 VSS.n16014 0.905
R18594 VSS.n16024 VSS.n16023 0.905
R18595 VSS.n16029 VSS.n16028 0.905
R18596 VSS.n15637 VSS.n15636 0.905
R18597 VSS.n15646 VSS.n15645 0.905
R18598 VSS.n15651 VSS.n15650 0.905
R18599 VSS.n15660 VSS.n15659 0.905
R18600 VSS.n15665 VSS.n15664 0.905
R18601 VSS.n15674 VSS.n15673 0.905
R18602 VSS.n15679 VSS.n15678 0.905
R18603 VSS.n15688 VSS.n15687 0.905
R18604 VSS.n15693 VSS.n15692 0.905
R18605 VSS.n15702 VSS.n15701 0.905
R18606 VSS.n15707 VSS.n15706 0.905
R18607 VSS.n15721 VSS.n15720 0.905
R18608 VSS.n15719 VSS.n14573 0.905
R18609 VSS.n14575 VSS.n14574 0.905
R18610 VSS.n14572 VSS.n14571 0.905
R18611 VSS.n15738 VSS.n15737 0.905
R18612 VSS.n15743 VSS.n15742 0.905
R18613 VSS.n15752 VSS.n15751 0.905
R18614 VSS.n15757 VSS.n15756 0.905
R18615 VSS.n15766 VSS.n15765 0.905
R18616 VSS.n15771 VSS.n15770 0.905
R18617 VSS.n15780 VSS.n15779 0.905
R18618 VSS.n15785 VSS.n15784 0.905
R18619 VSS.n15393 VSS.n15392 0.905
R18620 VSS.n15402 VSS.n15401 0.905
R18621 VSS.n15407 VSS.n15406 0.905
R18622 VSS.n15416 VSS.n15415 0.905
R18623 VSS.n15421 VSS.n15420 0.905
R18624 VSS.n15430 VSS.n15429 0.905
R18625 VSS.n15435 VSS.n15434 0.905
R18626 VSS.n15444 VSS.n15443 0.905
R18627 VSS.n15449 VSS.n15448 0.905
R18628 VSS.n15458 VSS.n15457 0.905
R18629 VSS.n15463 VSS.n15462 0.905
R18630 VSS.n15477 VSS.n15476 0.905
R18631 VSS.n15475 VSS.n14579 0.905
R18632 VSS.n14581 VSS.n14580 0.905
R18633 VSS.n14578 VSS.n14577 0.905
R18634 VSS.n15494 VSS.n15493 0.905
R18635 VSS.n15499 VSS.n15498 0.905
R18636 VSS.n15508 VSS.n15507 0.905
R18637 VSS.n15513 VSS.n15512 0.905
R18638 VSS.n15522 VSS.n15521 0.905
R18639 VSS.n15527 VSS.n15526 0.905
R18640 VSS.n15536 VSS.n15535 0.905
R18641 VSS.n15541 VSS.n15540 0.905
R18642 VSS.n15149 VSS.n15148 0.905
R18643 VSS.n15158 VSS.n15157 0.905
R18644 VSS.n15163 VSS.n15162 0.905
R18645 VSS.n15172 VSS.n15171 0.905
R18646 VSS.n15177 VSS.n15176 0.905
R18647 VSS.n15186 VSS.n15185 0.905
R18648 VSS.n15191 VSS.n15190 0.905
R18649 VSS.n15200 VSS.n15199 0.905
R18650 VSS.n15205 VSS.n15204 0.905
R18651 VSS.n15214 VSS.n15213 0.905
R18652 VSS.n15219 VSS.n15218 0.905
R18653 VSS.n15233 VSS.n15232 0.905
R18654 VSS.n15231 VSS.n14585 0.905
R18655 VSS.n14587 VSS.n14586 0.905
R18656 VSS.n14584 VSS.n14583 0.905
R18657 VSS.n15250 VSS.n15249 0.905
R18658 VSS.n15255 VSS.n15254 0.905
R18659 VSS.n15264 VSS.n15263 0.905
R18660 VSS.n15269 VSS.n15268 0.905
R18661 VSS.n15278 VSS.n15277 0.905
R18662 VSS.n15283 VSS.n15282 0.905
R18663 VSS.n15292 VSS.n15291 0.905
R18664 VSS.n15297 VSS.n15296 0.905
R18665 VSS.n14905 VSS.n14904 0.905
R18666 VSS.n14914 VSS.n14913 0.905
R18667 VSS.n14919 VSS.n14918 0.905
R18668 VSS.n14928 VSS.n14927 0.905
R18669 VSS.n14933 VSS.n14932 0.905
R18670 VSS.n14942 VSS.n14941 0.905
R18671 VSS.n14947 VSS.n14946 0.905
R18672 VSS.n14956 VSS.n14955 0.905
R18673 VSS.n14961 VSS.n14960 0.905
R18674 VSS.n14970 VSS.n14969 0.905
R18675 VSS.n14975 VSS.n14974 0.905
R18676 VSS.n14989 VSS.n14988 0.905
R18677 VSS.n14987 VSS.n14591 0.905
R18678 VSS.n14593 VSS.n14592 0.905
R18679 VSS.n14590 VSS.n14589 0.905
R18680 VSS.n15006 VSS.n15005 0.905
R18681 VSS.n15011 VSS.n15010 0.905
R18682 VSS.n15020 VSS.n15019 0.905
R18683 VSS.n15025 VSS.n15024 0.905
R18684 VSS.n15034 VSS.n15033 0.905
R18685 VSS.n15039 VSS.n15038 0.905
R18686 VSS.n15048 VSS.n15047 0.905
R18687 VSS.n15053 VSS.n15052 0.905
R18688 VSS.n14646 VSS.n14645 0.905
R18689 VSS.n14658 VSS.n14657 0.905
R18690 VSS.n14663 VSS.n14662 0.905
R18691 VSS.n14672 VSS.n14671 0.905
R18692 VSS.n14677 VSS.n14676 0.905
R18693 VSS.n14686 VSS.n14685 0.905
R18694 VSS.n14691 VSS.n14690 0.905
R18695 VSS.n14700 VSS.n14699 0.905
R18696 VSS.n14705 VSS.n14704 0.905
R18697 VSS.n14714 VSS.n14713 0.905
R18698 VSS.n14719 VSS.n14718 0.905
R18699 VSS.n14733 VSS.n14732 0.905
R18700 VSS.n14731 VSS.n14597 0.905
R18701 VSS.n14599 VSS.n14598 0.905
R18702 VSS.n14596 VSS.n14595 0.905
R18703 VSS.n14750 VSS.n14749 0.905
R18704 VSS.n14755 VSS.n14754 0.905
R18705 VSS.n14764 VSS.n14763 0.905
R18706 VSS.n14769 VSS.n14768 0.905
R18707 VSS.n14778 VSS.n14777 0.905
R18708 VSS.n14783 VSS.n14782 0.905
R18709 VSS.n14792 VSS.n14791 0.905
R18710 VSS.n14797 VSS.n14796 0.905
R18711 VSS.n12430 VSS.n12429 0.905
R18712 VSS.n12439 VSS.n12438 0.905
R18713 VSS.n12444 VSS.n12443 0.905
R18714 VSS.n12453 VSS.n12452 0.905
R18715 VSS.n12458 VSS.n12457 0.905
R18716 VSS.n12467 VSS.n12466 0.905
R18717 VSS.n12472 VSS.n12471 0.905
R18718 VSS.n12481 VSS.n12480 0.905
R18719 VSS.n12486 VSS.n12485 0.905
R18720 VSS.n12495 VSS.n12494 0.905
R18721 VSS.n12500 VSS.n12499 0.905
R18722 VSS.n12514 VSS.n12513 0.905
R18723 VSS.n12512 VSS.n10604 0.905
R18724 VSS.n10606 VSS.n10605 0.905
R18725 VSS.n10603 VSS.n10602 0.905
R18726 VSS.n12531 VSS.n12530 0.905
R18727 VSS.n12536 VSS.n12535 0.905
R18728 VSS.n12545 VSS.n12544 0.905
R18729 VSS.n12550 VSS.n12549 0.905
R18730 VSS.n12559 VSS.n12558 0.905
R18731 VSS.n12564 VSS.n12563 0.905
R18732 VSS.n12573 VSS.n12572 0.905
R18733 VSS.n12623 VSS.n12622 0.905
R18734 VSS.n12634 VSS.n12633 0.905
R18735 VSS.n12174 VSS.n12173 0.905
R18736 VSS.n12183 VSS.n12182 0.905
R18737 VSS.n12188 VSS.n12187 0.905
R18738 VSS.n12197 VSS.n12196 0.905
R18739 VSS.n12202 VSS.n12201 0.905
R18740 VSS.n12211 VSS.n12210 0.905
R18741 VSS.n12216 VSS.n12215 0.905
R18742 VSS.n12225 VSS.n12224 0.905
R18743 VSS.n12230 VSS.n12229 0.905
R18744 VSS.n12239 VSS.n12238 0.905
R18745 VSS.n12244 VSS.n12243 0.905
R18746 VSS.n12258 VSS.n12257 0.905
R18747 VSS.n12256 VSS.n10610 0.905
R18748 VSS.n10612 VSS.n10611 0.905
R18749 VSS.n10609 VSS.n10608 0.905
R18750 VSS.n12275 VSS.n12274 0.905
R18751 VSS.n12280 VSS.n12279 0.905
R18752 VSS.n12289 VSS.n12288 0.905
R18753 VSS.n12294 VSS.n12293 0.905
R18754 VSS.n12303 VSS.n12302 0.905
R18755 VSS.n12308 VSS.n12307 0.905
R18756 VSS.n12317 VSS.n12316 0.905
R18757 VSS.n12322 VSS.n12321 0.905
R18758 VSS.n11930 VSS.n11929 0.905
R18759 VSS.n11939 VSS.n11938 0.905
R18760 VSS.n11944 VSS.n11943 0.905
R18761 VSS.n11953 VSS.n11952 0.905
R18762 VSS.n11958 VSS.n11957 0.905
R18763 VSS.n11967 VSS.n11966 0.905
R18764 VSS.n11972 VSS.n11971 0.905
R18765 VSS.n11981 VSS.n11980 0.905
R18766 VSS.n11986 VSS.n11985 0.905
R18767 VSS.n11995 VSS.n11994 0.905
R18768 VSS.n12000 VSS.n11999 0.905
R18769 VSS.n12014 VSS.n12013 0.905
R18770 VSS.n12012 VSS.n10616 0.905
R18771 VSS.n10618 VSS.n10617 0.905
R18772 VSS.n10615 VSS.n10614 0.905
R18773 VSS.n12031 VSS.n12030 0.905
R18774 VSS.n12036 VSS.n12035 0.905
R18775 VSS.n12045 VSS.n12044 0.905
R18776 VSS.n12050 VSS.n12049 0.905
R18777 VSS.n12059 VSS.n12058 0.905
R18778 VSS.n12064 VSS.n12063 0.905
R18779 VSS.n12073 VSS.n12072 0.905
R18780 VSS.n12078 VSS.n12077 0.905
R18781 VSS.n11686 VSS.n11685 0.905
R18782 VSS.n11695 VSS.n11694 0.905
R18783 VSS.n11700 VSS.n11699 0.905
R18784 VSS.n11709 VSS.n11708 0.905
R18785 VSS.n11714 VSS.n11713 0.905
R18786 VSS.n11723 VSS.n11722 0.905
R18787 VSS.n11728 VSS.n11727 0.905
R18788 VSS.n11737 VSS.n11736 0.905
R18789 VSS.n11742 VSS.n11741 0.905
R18790 VSS.n11751 VSS.n11750 0.905
R18791 VSS.n11756 VSS.n11755 0.905
R18792 VSS.n11770 VSS.n11769 0.905
R18793 VSS.n11768 VSS.n10622 0.905
R18794 VSS.n10624 VSS.n10623 0.905
R18795 VSS.n10621 VSS.n10620 0.905
R18796 VSS.n11787 VSS.n11786 0.905
R18797 VSS.n11792 VSS.n11791 0.905
R18798 VSS.n11801 VSS.n11800 0.905
R18799 VSS.n11806 VSS.n11805 0.905
R18800 VSS.n11815 VSS.n11814 0.905
R18801 VSS.n11820 VSS.n11819 0.905
R18802 VSS.n11829 VSS.n11828 0.905
R18803 VSS.n11834 VSS.n11833 0.905
R18804 VSS.n11442 VSS.n11441 0.905
R18805 VSS.n11451 VSS.n11450 0.905
R18806 VSS.n11456 VSS.n11455 0.905
R18807 VSS.n11465 VSS.n11464 0.905
R18808 VSS.n11470 VSS.n11469 0.905
R18809 VSS.n11479 VSS.n11478 0.905
R18810 VSS.n11484 VSS.n11483 0.905
R18811 VSS.n11493 VSS.n11492 0.905
R18812 VSS.n11498 VSS.n11497 0.905
R18813 VSS.n11507 VSS.n11506 0.905
R18814 VSS.n11512 VSS.n11511 0.905
R18815 VSS.n11526 VSS.n11525 0.905
R18816 VSS.n11524 VSS.n10628 0.905
R18817 VSS.n10630 VSS.n10629 0.905
R18818 VSS.n10627 VSS.n10626 0.905
R18819 VSS.n11543 VSS.n11542 0.905
R18820 VSS.n11548 VSS.n11547 0.905
R18821 VSS.n11557 VSS.n11556 0.905
R18822 VSS.n11562 VSS.n11561 0.905
R18823 VSS.n11571 VSS.n11570 0.905
R18824 VSS.n11576 VSS.n11575 0.905
R18825 VSS.n11585 VSS.n11584 0.905
R18826 VSS.n11590 VSS.n11589 0.905
R18827 VSS.n11198 VSS.n11197 0.905
R18828 VSS.n11207 VSS.n11206 0.905
R18829 VSS.n11212 VSS.n11211 0.905
R18830 VSS.n11221 VSS.n11220 0.905
R18831 VSS.n11226 VSS.n11225 0.905
R18832 VSS.n11235 VSS.n11234 0.905
R18833 VSS.n11240 VSS.n11239 0.905
R18834 VSS.n11249 VSS.n11248 0.905
R18835 VSS.n11254 VSS.n11253 0.905
R18836 VSS.n11263 VSS.n11262 0.905
R18837 VSS.n11268 VSS.n11267 0.905
R18838 VSS.n11282 VSS.n11281 0.905
R18839 VSS.n11280 VSS.n10634 0.905
R18840 VSS.n10636 VSS.n10635 0.905
R18841 VSS.n10633 VSS.n10632 0.905
R18842 VSS.n11299 VSS.n11298 0.905
R18843 VSS.n11304 VSS.n11303 0.905
R18844 VSS.n11313 VSS.n11312 0.905
R18845 VSS.n11318 VSS.n11317 0.905
R18846 VSS.n11327 VSS.n11326 0.905
R18847 VSS.n11332 VSS.n11331 0.905
R18848 VSS.n11341 VSS.n11340 0.905
R18849 VSS.n11346 VSS.n11345 0.905
R18850 VSS.n10954 VSS.n10953 0.905
R18851 VSS.n10963 VSS.n10962 0.905
R18852 VSS.n10968 VSS.n10967 0.905
R18853 VSS.n10977 VSS.n10976 0.905
R18854 VSS.n10982 VSS.n10981 0.905
R18855 VSS.n10991 VSS.n10990 0.905
R18856 VSS.n10996 VSS.n10995 0.905
R18857 VSS.n11005 VSS.n11004 0.905
R18858 VSS.n11010 VSS.n11009 0.905
R18859 VSS.n11019 VSS.n11018 0.905
R18860 VSS.n11024 VSS.n11023 0.905
R18861 VSS.n11038 VSS.n11037 0.905
R18862 VSS.n11036 VSS.n10640 0.905
R18863 VSS.n10642 VSS.n10641 0.905
R18864 VSS.n10639 VSS.n10638 0.905
R18865 VSS.n11055 VSS.n11054 0.905
R18866 VSS.n11060 VSS.n11059 0.905
R18867 VSS.n11069 VSS.n11068 0.905
R18868 VSS.n11074 VSS.n11073 0.905
R18869 VSS.n11083 VSS.n11082 0.905
R18870 VSS.n11088 VSS.n11087 0.905
R18871 VSS.n11097 VSS.n11096 0.905
R18872 VSS.n11102 VSS.n11101 0.905
R18873 VSS.n10695 VSS.n10694 0.905
R18874 VSS.n10707 VSS.n10706 0.905
R18875 VSS.n10712 VSS.n10711 0.905
R18876 VSS.n10721 VSS.n10720 0.905
R18877 VSS.n10726 VSS.n10725 0.905
R18878 VSS.n10735 VSS.n10734 0.905
R18879 VSS.n10740 VSS.n10739 0.905
R18880 VSS.n10749 VSS.n10748 0.905
R18881 VSS.n10754 VSS.n10753 0.905
R18882 VSS.n10763 VSS.n10762 0.905
R18883 VSS.n10768 VSS.n10767 0.905
R18884 VSS.n10782 VSS.n10781 0.905
R18885 VSS.n10780 VSS.n10646 0.905
R18886 VSS.n10648 VSS.n10647 0.905
R18887 VSS.n10645 VSS.n10644 0.905
R18888 VSS.n10799 VSS.n10798 0.905
R18889 VSS.n10804 VSS.n10803 0.905
R18890 VSS.n10813 VSS.n10812 0.905
R18891 VSS.n10818 VSS.n10817 0.905
R18892 VSS.n10827 VSS.n10826 0.905
R18893 VSS.n10832 VSS.n10831 0.905
R18894 VSS.n10841 VSS.n10840 0.905
R18895 VSS.n10846 VSS.n10845 0.905
R18896 VSS.n8998 VSS.n8997 0.905
R18897 VSS.n9007 VSS.n9006 0.905
R18898 VSS.n9012 VSS.n9011 0.905
R18899 VSS.n9021 VSS.n9020 0.905
R18900 VSS.n9026 VSS.n9025 0.905
R18901 VSS.n9035 VSS.n9034 0.905
R18902 VSS.n9040 VSS.n9039 0.905
R18903 VSS.n9049 VSS.n9048 0.905
R18904 VSS.n9054 VSS.n9053 0.905
R18905 VSS.n9063 VSS.n9062 0.905
R18906 VSS.n9068 VSS.n9067 0.905
R18907 VSS.n9082 VSS.n9081 0.905
R18908 VSS.n9080 VSS.n7172 0.905
R18909 VSS.n7174 VSS.n7173 0.905
R18910 VSS.n7171 VSS.n7170 0.905
R18911 VSS.n9099 VSS.n9098 0.905
R18912 VSS.n9104 VSS.n9103 0.905
R18913 VSS.n9113 VSS.n9112 0.905
R18914 VSS.n9118 VSS.n9117 0.905
R18915 VSS.n9127 VSS.n9126 0.905
R18916 VSS.n9132 VSS.n9131 0.905
R18917 VSS.n9141 VSS.n9140 0.905
R18918 VSS.n9191 VSS.n9190 0.905
R18919 VSS.n9202 VSS.n9201 0.905
R18920 VSS.n8742 VSS.n8741 0.905
R18921 VSS.n8751 VSS.n8750 0.905
R18922 VSS.n8756 VSS.n8755 0.905
R18923 VSS.n8765 VSS.n8764 0.905
R18924 VSS.n8770 VSS.n8769 0.905
R18925 VSS.n8779 VSS.n8778 0.905
R18926 VSS.n8784 VSS.n8783 0.905
R18927 VSS.n8793 VSS.n8792 0.905
R18928 VSS.n8798 VSS.n8797 0.905
R18929 VSS.n8807 VSS.n8806 0.905
R18930 VSS.n8812 VSS.n8811 0.905
R18931 VSS.n8826 VSS.n8825 0.905
R18932 VSS.n8824 VSS.n7178 0.905
R18933 VSS.n7180 VSS.n7179 0.905
R18934 VSS.n7177 VSS.n7176 0.905
R18935 VSS.n8843 VSS.n8842 0.905
R18936 VSS.n8848 VSS.n8847 0.905
R18937 VSS.n8857 VSS.n8856 0.905
R18938 VSS.n8862 VSS.n8861 0.905
R18939 VSS.n8871 VSS.n8870 0.905
R18940 VSS.n8876 VSS.n8875 0.905
R18941 VSS.n8885 VSS.n8884 0.905
R18942 VSS.n8890 VSS.n8889 0.905
R18943 VSS.n8498 VSS.n8497 0.905
R18944 VSS.n8507 VSS.n8506 0.905
R18945 VSS.n8512 VSS.n8511 0.905
R18946 VSS.n8521 VSS.n8520 0.905
R18947 VSS.n8526 VSS.n8525 0.905
R18948 VSS.n8535 VSS.n8534 0.905
R18949 VSS.n8540 VSS.n8539 0.905
R18950 VSS.n8549 VSS.n8548 0.905
R18951 VSS.n8554 VSS.n8553 0.905
R18952 VSS.n8563 VSS.n8562 0.905
R18953 VSS.n8568 VSS.n8567 0.905
R18954 VSS.n8582 VSS.n8581 0.905
R18955 VSS.n8580 VSS.n7184 0.905
R18956 VSS.n7186 VSS.n7185 0.905
R18957 VSS.n7183 VSS.n7182 0.905
R18958 VSS.n8599 VSS.n8598 0.905
R18959 VSS.n8604 VSS.n8603 0.905
R18960 VSS.n8613 VSS.n8612 0.905
R18961 VSS.n8618 VSS.n8617 0.905
R18962 VSS.n8627 VSS.n8626 0.905
R18963 VSS.n8632 VSS.n8631 0.905
R18964 VSS.n8641 VSS.n8640 0.905
R18965 VSS.n8646 VSS.n8645 0.905
R18966 VSS.n8254 VSS.n8253 0.905
R18967 VSS.n8263 VSS.n8262 0.905
R18968 VSS.n8268 VSS.n8267 0.905
R18969 VSS.n8277 VSS.n8276 0.905
R18970 VSS.n8282 VSS.n8281 0.905
R18971 VSS.n8291 VSS.n8290 0.905
R18972 VSS.n8296 VSS.n8295 0.905
R18973 VSS.n8305 VSS.n8304 0.905
R18974 VSS.n8310 VSS.n8309 0.905
R18975 VSS.n8319 VSS.n8318 0.905
R18976 VSS.n8324 VSS.n8323 0.905
R18977 VSS.n8338 VSS.n8337 0.905
R18978 VSS.n8336 VSS.n7190 0.905
R18979 VSS.n7192 VSS.n7191 0.905
R18980 VSS.n7189 VSS.n7188 0.905
R18981 VSS.n8355 VSS.n8354 0.905
R18982 VSS.n8360 VSS.n8359 0.905
R18983 VSS.n8369 VSS.n8368 0.905
R18984 VSS.n8374 VSS.n8373 0.905
R18985 VSS.n8383 VSS.n8382 0.905
R18986 VSS.n8388 VSS.n8387 0.905
R18987 VSS.n8397 VSS.n8396 0.905
R18988 VSS.n8402 VSS.n8401 0.905
R18989 VSS.n8010 VSS.n8009 0.905
R18990 VSS.n8019 VSS.n8018 0.905
R18991 VSS.n8024 VSS.n8023 0.905
R18992 VSS.n8033 VSS.n8032 0.905
R18993 VSS.n8038 VSS.n8037 0.905
R18994 VSS.n8047 VSS.n8046 0.905
R18995 VSS.n8052 VSS.n8051 0.905
R18996 VSS.n8061 VSS.n8060 0.905
R18997 VSS.n8066 VSS.n8065 0.905
R18998 VSS.n8075 VSS.n8074 0.905
R18999 VSS.n8080 VSS.n8079 0.905
R19000 VSS.n8094 VSS.n8093 0.905
R19001 VSS.n8092 VSS.n7196 0.905
R19002 VSS.n7198 VSS.n7197 0.905
R19003 VSS.n7195 VSS.n7194 0.905
R19004 VSS.n8111 VSS.n8110 0.905
R19005 VSS.n8116 VSS.n8115 0.905
R19006 VSS.n8125 VSS.n8124 0.905
R19007 VSS.n8130 VSS.n8129 0.905
R19008 VSS.n8139 VSS.n8138 0.905
R19009 VSS.n8144 VSS.n8143 0.905
R19010 VSS.n8153 VSS.n8152 0.905
R19011 VSS.n8158 VSS.n8157 0.905
R19012 VSS.n7766 VSS.n7765 0.905
R19013 VSS.n7775 VSS.n7774 0.905
R19014 VSS.n7780 VSS.n7779 0.905
R19015 VSS.n7789 VSS.n7788 0.905
R19016 VSS.n7794 VSS.n7793 0.905
R19017 VSS.n7803 VSS.n7802 0.905
R19018 VSS.n7808 VSS.n7807 0.905
R19019 VSS.n7817 VSS.n7816 0.905
R19020 VSS.n7822 VSS.n7821 0.905
R19021 VSS.n7831 VSS.n7830 0.905
R19022 VSS.n7836 VSS.n7835 0.905
R19023 VSS.n7850 VSS.n7849 0.905
R19024 VSS.n7848 VSS.n7202 0.905
R19025 VSS.n7204 VSS.n7203 0.905
R19026 VSS.n7201 VSS.n7200 0.905
R19027 VSS.n7867 VSS.n7866 0.905
R19028 VSS.n7872 VSS.n7871 0.905
R19029 VSS.n7881 VSS.n7880 0.905
R19030 VSS.n7886 VSS.n7885 0.905
R19031 VSS.n7895 VSS.n7894 0.905
R19032 VSS.n7900 VSS.n7899 0.905
R19033 VSS.n7909 VSS.n7908 0.905
R19034 VSS.n7914 VSS.n7913 0.905
R19035 VSS.n7522 VSS.n7521 0.905
R19036 VSS.n7531 VSS.n7530 0.905
R19037 VSS.n7536 VSS.n7535 0.905
R19038 VSS.n7545 VSS.n7544 0.905
R19039 VSS.n7550 VSS.n7549 0.905
R19040 VSS.n7559 VSS.n7558 0.905
R19041 VSS.n7564 VSS.n7563 0.905
R19042 VSS.n7573 VSS.n7572 0.905
R19043 VSS.n7578 VSS.n7577 0.905
R19044 VSS.n7587 VSS.n7586 0.905
R19045 VSS.n7592 VSS.n7591 0.905
R19046 VSS.n7606 VSS.n7605 0.905
R19047 VSS.n7604 VSS.n7208 0.905
R19048 VSS.n7210 VSS.n7209 0.905
R19049 VSS.n7207 VSS.n7206 0.905
R19050 VSS.n7623 VSS.n7622 0.905
R19051 VSS.n7628 VSS.n7627 0.905
R19052 VSS.n7637 VSS.n7636 0.905
R19053 VSS.n7642 VSS.n7641 0.905
R19054 VSS.n7651 VSS.n7650 0.905
R19055 VSS.n7656 VSS.n7655 0.905
R19056 VSS.n7665 VSS.n7664 0.905
R19057 VSS.n7670 VSS.n7669 0.905
R19058 VSS.n7263 VSS.n7262 0.905
R19059 VSS.n7275 VSS.n7274 0.905
R19060 VSS.n7280 VSS.n7279 0.905
R19061 VSS.n7289 VSS.n7288 0.905
R19062 VSS.n7294 VSS.n7293 0.905
R19063 VSS.n7303 VSS.n7302 0.905
R19064 VSS.n7308 VSS.n7307 0.905
R19065 VSS.n7317 VSS.n7316 0.905
R19066 VSS.n7322 VSS.n7321 0.905
R19067 VSS.n7331 VSS.n7330 0.905
R19068 VSS.n7336 VSS.n7335 0.905
R19069 VSS.n7350 VSS.n7349 0.905
R19070 VSS.n7348 VSS.n7214 0.905
R19071 VSS.n7216 VSS.n7215 0.905
R19072 VSS.n7213 VSS.n7212 0.905
R19073 VSS.n7367 VSS.n7366 0.905
R19074 VSS.n7372 VSS.n7371 0.905
R19075 VSS.n7381 VSS.n7380 0.905
R19076 VSS.n7386 VSS.n7385 0.905
R19077 VSS.n7395 VSS.n7394 0.905
R19078 VSS.n7400 VSS.n7399 0.905
R19079 VSS.n7409 VSS.n7408 0.905
R19080 VSS.n7414 VSS.n7413 0.905
R19081 VSS.n1021 VSS.n1019 0.905
R19082 VSS.n1030 VSS.n1020 0.905
R19083 VSS.n1253 VSS.n1028 0.905
R19084 VSS.n1248 VSS.n1029 0.905
R19085 VSS.n1247 VSS.n1033 0.905
R19086 VSS.n1240 VSS.n1037 0.905
R19087 VSS.n1040 VSS.n1039 0.905
R19088 VSS.n1049 VSS.n1041 0.905
R19089 VSS.n1230 VSS.n1047 0.905
R19090 VSS.n1225 VSS.n1048 0.905
R19091 VSS.n1224 VSS.n1052 0.905
R19092 VSS.n1217 VSS.n1056 0.905
R19093 VSS.n1059 VSS.n1058 0.905
R19094 VSS.n1068 VSS.n1060 0.905
R19095 VSS.n1207 VSS.n1066 0.905
R19096 VSS.n1202 VSS.n1067 0.905
R19097 VSS.n1201 VSS.n1071 0.905
R19098 VSS.n1194 VSS.n1075 0.905
R19099 VSS.n1078 VSS.n1077 0.905
R19100 VSS.n1087 VSS.n1079 0.905
R19101 VSS.n1184 VSS.n1085 0.905
R19102 VSS.n1179 VSS.n1086 0.905
R19103 VSS.n1178 VSS.n1090 0.905
R19104 VSS.n1171 VSS.n1094 0.905
R19105 VSS.n921 VSS.n713 0.905
R19106 VSS.n926 VSS.n711 0.905
R19107 VSS.n927 VSS.n706 0.905
R19108 VSS.n935 VSS.n934 0.905
R19109 VSS.n939 VSS.n704 0.905
R19110 VSS.n946 VSS.n700 0.905
R19111 VSS.n945 VSS.n696 0.905
R19112 VSS.n698 VSS.n697 0.905
R19113 VSS.n956 VSS.n692 0.905
R19114 VSS.n961 VSS.n690 0.905
R19115 VSS.n962 VSS.n685 0.905
R19116 VSS.n970 VSS.n969 0.905
R19117 VSS.n974 VSS.n683 0.905
R19118 VSS.n981 VSS.n679 0.905
R19119 VSS.n980 VSS.n675 0.905
R19120 VSS.n677 VSS.n676 0.905
R19121 VSS.n991 VSS.n671 0.905
R19122 VSS.n996 VSS.n669 0.905
R19123 VSS.n997 VSS.n664 0.905
R19124 VSS.n1005 VSS.n1004 0.905
R19125 VSS.n1009 VSS.n662 0.905
R19126 VSS.n1016 VSS.n658 0.905
R19127 VSS.n1015 VSS.n655 0.905
R19128 VSS.n1262 VSS.n656 0.905
R19129 VSS.n778 VSS.n590 0.905
R19130 VSS.n788 VSS.n787 0.905
R19131 VSS.n792 VSS.n776 0.905
R19132 VSS.n799 VSS.n772 0.905
R19133 VSS.n798 VSS.n768 0.905
R19134 VSS.n770 VSS.n769 0.905
R19135 VSS.n809 VSS.n764 0.905
R19136 VSS.n814 VSS.n762 0.905
R19137 VSS.n815 VSS.n757 0.905
R19138 VSS.n823 VSS.n822 0.905
R19139 VSS.n827 VSS.n755 0.905
R19140 VSS.n834 VSS.n751 0.905
R19141 VSS.n833 VSS.n747 0.905
R19142 VSS.n749 VSS.n748 0.905
R19143 VSS.n844 VSS.n743 0.905
R19144 VSS.n849 VSS.n741 0.905
R19145 VSS.n850 VSS.n736 0.905
R19146 VSS.n858 VSS.n857 0.905
R19147 VSS.n862 VSS.n734 0.905
R19148 VSS.n869 VSS.n730 0.905
R19149 VSS.n868 VSS.n725 0.905
R19150 VSS.n728 VSS.n727 0.905
R19151 VSS.n726 VSS.n721 0.905
R19152 VSS.n884 VSS.n719 0.905
R19153 VSS.n5605 VSS.n1380 0.905
R19154 VSS.n5601 VSS.n5600 0.905
R19155 VSS.n5599 VSS.n521 0.905
R19156 VSS.n530 VSS.n522 0.905
R19157 VSS.n5776 VSS.n528 0.905
R19158 VSS.n5771 VSS.n529 0.905
R19159 VSS.n5770 VSS.n533 0.905
R19160 VSS.n5763 VSS.n537 0.905
R19161 VSS.n540 VSS.n539 0.905
R19162 VSS.n549 VSS.n541 0.905
R19163 VSS.n5753 VSS.n547 0.905
R19164 VSS.n5748 VSS.n548 0.905
R19165 VSS.n5747 VSS.n552 0.905
R19166 VSS.n5740 VSS.n556 0.905
R19167 VSS.n559 VSS.n558 0.905
R19168 VSS.n568 VSS.n560 0.905
R19169 VSS.n5730 VSS.n566 0.905
R19170 VSS.n5725 VSS.n567 0.905
R19171 VSS.n5724 VSS.n571 0.905
R19172 VSS.n5717 VSS.n575 0.905
R19173 VSS.n578 VSS.n577 0.905
R19174 VSS.n587 VSS.n579 0.905
R19175 VSS.n5707 VSS.n585 0.905
R19176 VSS.n5702 VSS.n586 0.905
R19177 VSS.n5494 VSS.n1441 0.905
R19178 VSS.n5502 VSS.n5501 0.905
R19179 VSS.n5506 VSS.n1439 0.905
R19180 VSS.n5513 VSS.n1435 0.905
R19181 VSS.n5512 VSS.n1431 0.905
R19182 VSS.n1433 VSS.n1432 0.905
R19183 VSS.n5523 VSS.n1427 0.905
R19184 VSS.n5528 VSS.n1425 0.905
R19185 VSS.n5529 VSS.n1420 0.905
R19186 VSS.n5537 VSS.n5536 0.905
R19187 VSS.n5541 VSS.n1418 0.905
R19188 VSS.n5548 VSS.n1414 0.905
R19189 VSS.n5547 VSS.n1410 0.905
R19190 VSS.n1412 VSS.n1411 0.905
R19191 VSS.n5558 VSS.n1406 0.905
R19192 VSS.n5563 VSS.n1404 0.905
R19193 VSS.n5564 VSS.n1399 0.905
R19194 VSS.n5572 VSS.n5571 0.905
R19195 VSS.n5576 VSS.n1397 0.905
R19196 VSS.n5584 VSS.n1391 0.905
R19197 VSS.n5583 VSS.n1392 0.905
R19198 VSS.n5589 VSS.n5588 0.905
R19199 VSS.n5590 VSS.n1384 0.905
R19200 VSS.n5616 VSS.n1382 0.905
R19201 VSS.n5397 VSS.n1521 0.905
R19202 VSS.n5392 VSS.n5237 0.905
R19203 VSS.n5391 VSS.n5239 0.905
R19204 VSS.n5384 VSS.n5244 0.905
R19205 VSS.n5247 VSS.n5246 0.905
R19206 VSS.n5256 VSS.n5248 0.905
R19207 VSS.n5374 VSS.n5254 0.905
R19208 VSS.n5369 VSS.n5255 0.905
R19209 VSS.n5368 VSS.n5259 0.905
R19210 VSS.n5361 VSS.n5263 0.905
R19211 VSS.n5266 VSS.n5265 0.905
R19212 VSS.n5275 VSS.n5267 0.905
R19213 VSS.n5351 VSS.n5273 0.905
R19214 VSS.n5346 VSS.n5274 0.905
R19215 VSS.n5345 VSS.n5278 0.905
R19216 VSS.n5338 VSS.n5282 0.905
R19217 VSS.n5285 VSS.n5284 0.905
R19218 VSS.n5294 VSS.n5286 0.905
R19219 VSS.n5328 VSS.n5292 0.905
R19220 VSS.n5323 VSS.n5293 0.905
R19221 VSS.n5322 VSS.n5297 0.905
R19222 VSS.n5315 VSS.n5301 0.905
R19223 VSS.n5305 VSS.n5304 0.905
R19224 VSS.n5306 VSS.n1446 0.905
R19225 VSS.n5135 VSS.n1582 0.905
R19226 VSS.n5143 VSS.n5142 0.905
R19227 VSS.n5147 VSS.n1580 0.905
R19228 VSS.n5154 VSS.n1576 0.905
R19229 VSS.n5153 VSS.n1572 0.905
R19230 VSS.n1574 VSS.n1573 0.905
R19231 VSS.n5164 VSS.n1568 0.905
R19232 VSS.n5169 VSS.n1566 0.905
R19233 VSS.n5170 VSS.n1561 0.905
R19234 VSS.n5178 VSS.n5177 0.905
R19235 VSS.n5182 VSS.n1559 0.905
R19236 VSS.n5189 VSS.n1555 0.905
R19237 VSS.n5188 VSS.n1551 0.905
R19238 VSS.n1553 VSS.n1552 0.905
R19239 VSS.n5199 VSS.n1547 0.905
R19240 VSS.n5204 VSS.n1545 0.905
R19241 VSS.n5205 VSS.n1540 0.905
R19242 VSS.n5213 VSS.n5212 0.905
R19243 VSS.n5217 VSS.n1538 0.905
R19244 VSS.n5225 VSS.n1532 0.905
R19245 VSS.n5224 VSS.n1533 0.905
R19246 VSS.n5230 VSS.n5229 0.905
R19247 VSS.n5231 VSS.n1525 0.905
R19248 VSS.n5408 VSS.n1523 0.905
R19249 VSS.n4766 VSS.n4762 0.905
R19250 VSS.n4774 VSS.n4763 0.905
R19251 VSS.n4920 VSS.n4772 0.905
R19252 VSS.n4915 VSS.n4773 0.905
R19253 VSS.n4914 VSS.n4777 0.905
R19254 VSS.n4907 VSS.n4781 0.905
R19255 VSS.n4784 VSS.n4783 0.905
R19256 VSS.n4793 VSS.n4785 0.905
R19257 VSS.n4897 VSS.n4791 0.905
R19258 VSS.n4892 VSS.n4792 0.905
R19259 VSS.n4891 VSS.n4796 0.905
R19260 VSS.n4884 VSS.n4800 0.905
R19261 VSS.n4803 VSS.n4802 0.905
R19262 VSS.n4812 VSS.n4804 0.905
R19263 VSS.n4874 VSS.n4810 0.905
R19264 VSS.n4869 VSS.n4811 0.905
R19265 VSS.n4868 VSS.n4815 0.905
R19266 VSS.n4861 VSS.n4819 0.905
R19267 VSS.n4822 VSS.n4821 0.905
R19268 VSS.n4831 VSS.n4823 0.905
R19269 VSS.n4851 VSS.n4829 0.905
R19270 VSS.n4846 VSS.n4830 0.905
R19271 VSS.n4845 VSS.n4834 0.905
R19272 VSS.n4838 VSS.n4836 0.905
R19273 VSS.n4651 VSS.n3155 0.905
R19274 VSS.n4662 VSS.n4652 0.905
R19275 VSS.n5013 VSS.n4660 0.905
R19276 VSS.n5008 VSS.n4661 0.905
R19277 VSS.n5007 VSS.n4665 0.905
R19278 VSS.n5000 VSS.n4669 0.905
R19279 VSS.n4672 VSS.n4671 0.905
R19280 VSS.n4681 VSS.n4673 0.905
R19281 VSS.n4990 VSS.n4679 0.905
R19282 VSS.n4985 VSS.n4680 0.905
R19283 VSS.n4984 VSS.n4684 0.905
R19284 VSS.n4977 VSS.n4688 0.905
R19285 VSS.n4691 VSS.n4690 0.905
R19286 VSS.n4700 VSS.n4692 0.905
R19287 VSS.n4967 VSS.n4698 0.905
R19288 VSS.n4962 VSS.n4699 0.905
R19289 VSS.n4961 VSS.n4703 0.905
R19290 VSS.n4954 VSS.n4707 0.905
R19291 VSS.n4710 VSS.n4709 0.905
R19292 VSS.n4719 VSS.n4711 0.905
R19293 VSS.n4944 VSS.n4717 0.905
R19294 VSS.n4939 VSS.n4718 0.905
R19295 VSS.n4938 VSS.n4722 0.905
R19296 VSS.n4931 VSS.n4726 0.905
R19297 VSS.n4547 VSS.n3218 0.905
R19298 VSS.n4554 VSS.n3214 0.905
R19299 VSS.n4553 VSS.n3210 0.905
R19300 VSS.n3212 VSS.n3211 0.905
R19301 VSS.n4564 VSS.n3206 0.905
R19302 VSS.n4569 VSS.n3204 0.905
R19303 VSS.n4570 VSS.n3199 0.905
R19304 VSS.n4578 VSS.n4577 0.905
R19305 VSS.n4582 VSS.n3197 0.905
R19306 VSS.n4589 VSS.n3193 0.905
R19307 VSS.n4588 VSS.n3189 0.905
R19308 VSS.n3191 VSS.n3190 0.905
R19309 VSS.n4599 VSS.n3185 0.905
R19310 VSS.n4604 VSS.n3183 0.905
R19311 VSS.n4605 VSS.n3178 0.905
R19312 VSS.n4613 VSS.n4612 0.905
R19313 VSS.n4617 VSS.n3176 0.905
R19314 VSS.n4624 VSS.n3172 0.905
R19315 VSS.n4623 VSS.n3168 0.905
R19316 VSS.n3170 VSS.n3169 0.905
R19317 VSS.n4634 VSS.n3164 0.905
R19318 VSS.n4639 VSS.n3162 0.905
R19319 VSS.n4640 VSS.n3158 0.905
R19320 VSS.n4647 VSS.n3156 0.905
R19321 VSS.n4176 VSS.n4172 0.905
R19322 VSS.n4184 VSS.n4173 0.905
R19323 VSS.n4311 VSS.n4182 0.905
R19324 VSS.n4306 VSS.n4183 0.905
R19325 VSS.n4305 VSS.n4187 0.905
R19326 VSS.n4298 VSS.n4191 0.905
R19327 VSS.n4194 VSS.n4193 0.905
R19328 VSS.n4203 VSS.n4195 0.905
R19329 VSS.n4288 VSS.n4201 0.905
R19330 VSS.n4283 VSS.n4202 0.905
R19331 VSS.n4282 VSS.n4206 0.905
R19332 VSS.n4275 VSS.n4210 0.905
R19333 VSS.n4213 VSS.n4212 0.905
R19334 VSS.n4222 VSS.n4214 0.905
R19335 VSS.n4265 VSS.n4220 0.905
R19336 VSS.n4260 VSS.n4221 0.905
R19337 VSS.n4259 VSS.n4225 0.905
R19338 VSS.n4252 VSS.n4229 0.905
R19339 VSS.n4232 VSS.n4231 0.905
R19340 VSS.n4238 VSS.n4233 0.905
R19341 VSS.n4242 VSS.n4237 0.905
R19342 VSS.n4537 VSS.n3223 0.905
R19343 VSS.n4536 VSS.n3224 0.905
R19344 VSS.n4542 VSS.n4541 0.905
R19345 VSS.n4063 VSS.n4061 0.905
R19346 VSS.n4072 VSS.n4062 0.905
R19347 VSS.n4404 VSS.n4070 0.905
R19348 VSS.n4399 VSS.n4071 0.905
R19349 VSS.n4398 VSS.n4075 0.905
R19350 VSS.n4391 VSS.n4079 0.905
R19351 VSS.n4082 VSS.n4081 0.905
R19352 VSS.n4091 VSS.n4083 0.905
R19353 VSS.n4381 VSS.n4089 0.905
R19354 VSS.n4376 VSS.n4090 0.905
R19355 VSS.n4375 VSS.n4094 0.905
R19356 VSS.n4368 VSS.n4098 0.905
R19357 VSS.n4101 VSS.n4100 0.905
R19358 VSS.n4110 VSS.n4102 0.905
R19359 VSS.n4358 VSS.n4108 0.905
R19360 VSS.n4353 VSS.n4109 0.905
R19361 VSS.n4352 VSS.n4113 0.905
R19362 VSS.n4345 VSS.n4117 0.905
R19363 VSS.n4120 VSS.n4119 0.905
R19364 VSS.n4129 VSS.n4121 0.905
R19365 VSS.n4335 VSS.n4127 0.905
R19366 VSS.n4330 VSS.n4128 0.905
R19367 VSS.n4329 VSS.n4132 0.905
R19368 VSS.n4322 VSS.n4136 0.905
R19369 VSS.n3963 VSS.n3383 0.905
R19370 VSS.n3968 VSS.n3381 0.905
R19371 VSS.n3969 VSS.n3376 0.905
R19372 VSS.n3977 VSS.n3976 0.905
R19373 VSS.n3981 VSS.n3374 0.905
R19374 VSS.n3988 VSS.n3370 0.905
R19375 VSS.n3987 VSS.n3366 0.905
R19376 VSS.n3368 VSS.n3367 0.905
R19377 VSS.n3998 VSS.n3362 0.905
R19378 VSS.n4003 VSS.n3360 0.905
R19379 VSS.n4004 VSS.n3355 0.905
R19380 VSS.n4012 VSS.n4011 0.905
R19381 VSS.n4016 VSS.n3353 0.905
R19382 VSS.n4023 VSS.n3349 0.905
R19383 VSS.n4022 VSS.n3345 0.905
R19384 VSS.n3347 VSS.n3346 0.905
R19385 VSS.n4033 VSS.n3341 0.905
R19386 VSS.n4038 VSS.n3339 0.905
R19387 VSS.n4039 VSS.n3334 0.905
R19388 VSS.n4047 VSS.n4046 0.905
R19389 VSS.n4051 VSS.n3332 0.905
R19390 VSS.n4058 VSS.n3328 0.905
R19391 VSS.n4057 VSS.n3325 0.905
R19392 VSS.n4413 VSS.n3326 0.905
R19393 VSS.n3564 VSS.n3560 0.905
R19394 VSS.n3572 VSS.n3561 0.905
R19395 VSS.n3707 VSS.n3570 0.905
R19396 VSS.n3702 VSS.n3571 0.905
R19397 VSS.n3701 VSS.n3575 0.905
R19398 VSS.n3694 VSS.n3579 0.905
R19399 VSS.n3582 VSS.n3581 0.905
R19400 VSS.n3591 VSS.n3583 0.905
R19401 VSS.n3684 VSS.n3589 0.905
R19402 VSS.n3679 VSS.n3590 0.905
R19403 VSS.n3678 VSS.n3594 0.905
R19404 VSS.n3671 VSS.n3598 0.905
R19405 VSS.n3601 VSS.n3600 0.905
R19406 VSS.n3610 VSS.n3602 0.905
R19407 VSS.n3661 VSS.n3608 0.905
R19408 VSS.n3656 VSS.n3609 0.905
R19409 VSS.n3655 VSS.n3613 0.905
R19410 VSS.n3648 VSS.n3617 0.905
R19411 VSS.n3620 VSS.n3619 0.905
R19412 VSS.n3633 VSS.n3621 0.905
R19413 VSS.n3638 VSS.n3627 0.905
R19414 VSS.n3632 VSS.n3631 0.905
R19415 VSS.n3630 VSS.n3389 0.905
R19416 VSS.n3952 VSS.n3390 0.905
R19417 VSS.n3808 VSS.n3807 0.905
R19418 VSS.n3460 VSS.n3452 0.905
R19419 VSS.n3800 VSS.n3457 0.905
R19420 VSS.n3795 VSS.n3458 0.905
R19421 VSS.n3794 VSS.n3463 0.905
R19422 VSS.n3787 VSS.n3467 0.905
R19423 VSS.n3470 VSS.n3469 0.905
R19424 VSS.n3479 VSS.n3471 0.905
R19425 VSS.n3777 VSS.n3477 0.905
R19426 VSS.n3772 VSS.n3478 0.905
R19427 VSS.n3771 VSS.n3482 0.905
R19428 VSS.n3764 VSS.n3486 0.905
R19429 VSS.n3489 VSS.n3488 0.905
R19430 VSS.n3498 VSS.n3490 0.905
R19431 VSS.n3754 VSS.n3496 0.905
R19432 VSS.n3749 VSS.n3497 0.905
R19433 VSS.n3748 VSS.n3501 0.905
R19434 VSS.n3741 VSS.n3505 0.905
R19435 VSS.n3508 VSS.n3507 0.905
R19436 VSS.n3517 VSS.n3509 0.905
R19437 VSS.n3731 VSS.n3515 0.905
R19438 VSS.n3726 VSS.n3516 0.905
R19439 VSS.n3725 VSS.n3520 0.905
R19440 VSS.n3718 VSS.n3524 0.905
R19441 VSS.n17768 VSS.n17767 0.855
R19442 VSS.n18103 VSS.n18102 0.852
R19443 VSS.n18103 VSS.n18098 0.852
R19444 VSS.n18103 VSS.n24 0.852
R19445 VSS.n18103 VSS.n26 0.852
R19446 VSS.n18103 VSS.n29 0.852
R19447 VSS.n18103 VSS.n18096 0.852
R19448 VSS.n17658 VSS.n17657 0.852
R19449 VSS.n17658 VSS.n17653 0.852
R19450 VSS.n17658 VSS.n17624 0.852
R19451 VSS.n17658 VSS.n17626 0.852
R19452 VSS.n17658 VSS.n17629 0.852
R19453 VSS.n17658 VSS.n17649 0.852
R19454 VSS.n17669 VSS.n17668 0.852
R19455 VSS.n17669 VSS.n17663 0.852
R19456 VSS.n17669 VSS.n14114 0.852
R19457 VSS.n17669 VSS.n14116 0.852
R19458 VSS.n17669 VSS.n14118 0.852
R19459 VSS.n17669 VSS.n17617 0.852
R19460 VSS.n17679 VSS.n17678 0.852
R19461 VSS.n17679 VSS.n17674 0.852
R19462 VSS.n17679 VSS.n10592 0.852
R19463 VSS.n17679 VSS.n10594 0.852
R19464 VSS.n17679 VSS.n10597 0.852
R19465 VSS.n17679 VSS.n14107 0.852
R19466 VSS.n17690 VSS.n17689 0.852
R19467 VSS.n17690 VSS.n17684 0.852
R19468 VSS.n17690 VSS.n7074 0.852
R19469 VSS.n17690 VSS.n7076 0.852
R19470 VSS.n17690 VSS.n7078 0.852
R19471 VSS.n17690 VSS.n10585 0.852
R19472 VSS.n17701 VSS.n17700 0.852
R19473 VSS.n17701 VSS.n17695 0.852
R19474 VSS.n17701 VSS.n511 0.852
R19475 VSS.n17701 VSS.n513 0.852
R19476 VSS.n17701 VSS.n515 0.852
R19477 VSS.n17701 VSS.n7067 0.852
R19478 VSS.n17712 VSS.n17711 0.852
R19479 VSS.n17712 VSS.n17706 0.852
R19480 VSS.n17712 VSS.n453 0.852
R19481 VSS.n17712 VSS.n455 0.852
R19482 VSS.n17712 VSS.n457 0.852
R19483 VSS.n17712 VSS.n504 0.852
R19484 VSS.n17722 VSS.n17721 0.852
R19485 VSS.n17722 VSS.n17717 0.852
R19486 VSS.n17722 VSS.n314 0.852
R19487 VSS.n17722 VSS.n316 0.852
R19488 VSS.n17722 VSS.n319 0.852
R19489 VSS.n17722 VSS.n446 0.852
R19490 VSS.n17733 VSS.n17732 0.852
R19491 VSS.n17733 VSS.n17727 0.852
R19492 VSS.n17733 VSS.n303 0.852
R19493 VSS.n17733 VSS.n307 0.852
R19494 VSS.n17734 VSS.n17733 0.852
R19495 VSS.n18103 VSS.n18100 0.849
R19496 VSS.n17658 VSS.n17655 0.849
R19497 VSS.n17669 VSS.n17666 0.849
R19498 VSS.n17679 VSS.n17676 0.849
R19499 VSS.n17690 VSS.n17687 0.849
R19500 VSS.n17701 VSS.n17698 0.849
R19501 VSS.n17712 VSS.n17709 0.849
R19502 VSS.n17722 VSS.n17719 0.849
R19503 VSS.n17733 VSS.n305 0.849
R19504 VSS.n17733 VSS.n17730 0.849
R19505 VSS.n18324 VSS.n18323 0.849
R19506 VSS.n18324 VSS.n18315 0.849
R19507 VSS.n18324 VSS.n18313 0.849
R19508 VSS.n18324 VSS.n18310 0.849
R19509 VSS.n18324 VSS.n18308 0.849
R19510 VSS.n18324 VSS.n18305 0.849
R19511 VSS.n18324 VSS.n18303 0.849
R19512 VSS.n240 VSS.n222 0.849
R19513 VSS.n240 VSS.n226 0.849
R19514 VSS.n240 VSS.n215 0.849
R19515 VSS.n240 VSS.n229 0.849
R19516 VSS.n240 VSS.n213 0.849
R19517 VSS.n240 VSS.n232 0.849
R19518 VSS.n240 VSS.n210 0.849
R19519 VSS.n240 VSS.n239 0.849
R19520 VSS.n18258 VSS.n18257 0.849
R19521 VSS.n18258 VSS.n18248 0.849
R19522 VSS.n18258 VSS.n18246 0.849
R19523 VSS.n18258 VSS.n18243 0.849
R19524 VSS.n18258 VSS.n18241 0.849
R19525 VSS.n18258 VSS.n18238 0.849
R19526 VSS.n18258 VSS.n18236 0.849
R19527 VSS.n14312 VSS.n14299 0.785
R19528 VSS.n17430 VSS.n17429 0.785
R19529 VSS.n17262 VSS.n17261 0.785
R19530 VSS.n17094 VSS.n17093 0.785
R19531 VSS.n16926 VSS.n16925 0.785
R19532 VSS.n16758 VSS.n16757 0.785
R19533 VSS.n12829 VSS.n12816 0.785
R19534 VSS.n13009 VSS.n12996 0.785
R19535 VSS.n13189 VSS.n13176 0.785
R19536 VSS.n13369 VSS.n13356 0.785
R19537 VSS.n13549 VSS.n13536 0.785
R19538 VSS.n13729 VSS.n13716 0.785
R19539 VSS.n13909 VSS.n13896 0.785
R19540 VSS.n10395 VSS.n10382 0.785
R19541 VSS.n10228 VSS.n10214 0.785
R19542 VSS.n10060 VSS.n10046 0.785
R19543 VSS.n9892 VSS.n9878 0.785
R19544 VSS.n9724 VSS.n9710 0.785
R19545 VSS.n9556 VSS.n9542 0.785
R19546 VSS.n9388 VSS.n9374 0.785
R19547 VSS.n2464 VSS.n2463 0.785
R19548 VSS.n2554 VSS.n2553 0.785
R19549 VSS.n2644 VSS.n2643 0.785
R19550 VSS.n2734 VSS.n2733 0.785
R19551 VSS.n2824 VSS.n2823 0.785
R19552 VSS.n2914 VSS.n2913 0.785
R19553 VSS.n3004 VSS.n3003 0.785
R19554 VSS.n6758 VSS.n6757 0.785
R19555 VSS.n6848 VSS.n6847 0.785
R19556 VSS.n6381 VSS.n6380 0.785
R19557 VSS.n6317 VSS.n6316 0.785
R19558 VSS.n6253 VSS.n6252 0.785
R19559 VSS.n6938 VSS.n6937 0.784
R19560 VSS.n402 VSS.n401 0.752
R19561 VSS.n403 VSS.n402 0.752
R19562 VSS.n411 VSS.n358 0.752
R19563 VSS.n411 VSS.n356 0.752
R19564 VSS.n18194 VSS.n18193 0.752
R19565 VSS.n18195 VSS.n18194 0.752
R19566 VSS.n18203 VSS.n18150 0.752
R19567 VSS.n18203 VSS.n18148 0.752
R19568 VSS VSS.n18025 0.737
R19569 VSS.n14460 VSS.n14459 0.735
R19570 VSS.n14280 VSS.n14279 0.735
R19571 VSS.n14057 VSS.n14056 0.735
R19572 VSS.n13877 VSS.n13876 0.735
R19573 VSS.n13697 VSS.n13696 0.735
R19574 VSS.n13517 VSS.n13516 0.735
R19575 VSS.n13337 VSS.n13336 0.735
R19576 VSS.n13157 VSS.n13156 0.735
R19577 VSS.n12977 VSS.n12976 0.735
R19578 VSS.n12797 VSS.n12796 0.735
R19579 VSS.n9227 VSS.n9226 0.735
R19580 VSS.n9395 VSS.n9394 0.735
R19581 VSS.n9563 VSS.n9562 0.735
R19582 VSS.n9731 VSS.n9730 0.735
R19583 VSS.n9899 VSS.n9898 0.735
R19584 VSS.n10067 VSS.n10066 0.735
R19585 VSS.n10235 VSS.n10234 0.735
R19586 VSS.n6931 VSS.n6402 0.735
R19587 VSS.n6841 VSS.n6492 0.735
R19588 VSS.n6751 VSS.n6582 0.735
R19589 VSS.n18042 VSS.n18041 0.677
R19590 VSS.n18127 VSS.n18110 0.677
R19591 VSS.n17598 VSS.n14479 0.569
R19592 VSS.n18047 VSS.n206 0.563
R19593 VSS.n18047 VSS.n204 0.563
R19594 VSS.n18047 VSS.n198 0.563
R19595 VSS.n18052 VSS.n185 0.563
R19596 VSS.n18052 VSS.n183 0.563
R19597 VSS.n18052 VSS.n177 0.563
R19598 VSS.n18057 VSS.n164 0.563
R19599 VSS.n18057 VSS.n162 0.563
R19600 VSS.n18057 VSS.n156 0.563
R19601 VSS.n18062 VSS.n143 0.563
R19602 VSS.n18062 VSS.n141 0.563
R19603 VSS.n18062 VSS.n135 0.563
R19604 VSS.n18067 VSS.n122 0.563
R19605 VSS.n18067 VSS.n120 0.563
R19606 VSS.n18067 VSS.n114 0.563
R19607 VSS.n18072 VSS.n101 0.563
R19608 VSS.n18072 VSS.n99 0.563
R19609 VSS.n18072 VSS.n93 0.563
R19610 VSS.n18077 VSS.n80 0.563
R19611 VSS.n18077 VSS.n78 0.563
R19612 VSS.n18077 VSS.n72 0.563
R19613 VSS.n18084 VSS.n18082 0.563
R19614 VSS.n18082 VSS.n59 0.563
R19615 VSS.n18082 VSS.n53 0.563
R19616 VSS.n292 VSS.n275 0.563
R19617 VSS.n292 VSS.n280 0.563
R19618 VSS.n292 VSS.n291 0.563
R19619 VSS.n18285 VSS.n18274 0.563
R19620 VSS.n18285 VSS.n18279 0.563
R19621 VSS.n18285 VSS.n18284 0.563
R19622 VSS.n18287 VSS.n18285 0.563
R19623 VSS.n14382 VSS 0.533
R19624 VSS.n14202 VSS 0.533
R19625 VSS VSS.n17472 0.533
R19626 VSS VSS.n17304 0.533
R19627 VSS VSS.n17136 0.533
R19628 VSS VSS.n16968 0.533
R19629 VSS VSS.n16800 0.533
R19630 VSS VSS.n16632 0.533
R19631 VSS.n13979 VSS 0.533
R19632 VSS.n13799 VSS 0.533
R19633 VSS.n13619 VSS 0.533
R19634 VSS.n13439 VSS 0.533
R19635 VSS.n13259 VSS 0.533
R19636 VSS.n13079 VSS 0.533
R19637 VSS.n12899 VSS 0.533
R19638 VSS.n12719 VSS 0.533
R19639 VSS VSS.n9262 0.533
R19640 VSS VSS.n9430 0.533
R19641 VSS VSS.n9598 0.533
R19642 VSS VSS.n9766 0.533
R19643 VSS VSS.n9934 0.533
R19644 VSS VSS.n10102 0.533
R19645 VSS VSS.n10270 0.533
R19646 VSS VSS.n10437 0.533
R19647 VSS VSS.n2424 0.533
R19648 VSS VSS.n2514 0.533
R19649 VSS VSS.n2604 0.533
R19650 VSS VSS.n2694 0.533
R19651 VSS VSS.n2784 0.533
R19652 VSS VSS.n2874 0.533
R19653 VSS VSS.n2964 0.533
R19654 VSS VSS.n3054 0.533
R19655 VSS.n6168 VSS 0.533
R19656 VSS.n6052 VSS 0.533
R19657 VSS.n5936 VSS 0.533
R19658 VSS.n5821 VSS 0.533
R19659 VSS VSS.n6897 0.533
R19660 VSS VSS.n6807 0.533
R19661 VSS VSS.n6717 0.533
R19662 VSS.n18019 VSS.n17923 0.533
R19663 VSS.n438 VSS 0.522
R19664 VSS.n494 VSS.n471 0.407
R19665 VSS.n18231 VSS 0.389
R19666 VSS VSS.n7060 0.385
R19667 VSS.n5132 VSS.n5131 0.366
R19668 VSS.n16589 VSS.n16588 0.357
R19669 VSS.n14081 VSS.n12637 0.357
R19670 VSS.n9206 VSS.n9205 0.357
R19671 VSS.n7046 VSS.n5784 0.357
R19672 VSS.n17754 VSS.n17753 0.352
R19673 VSS.n18022 VSS.n18021 0.348
R19674 VSS.n7060 VSS 0.331
R19675 VSS.n18231 VSS 0.331
R19676 VSS.n18026 VSS 0.33
R19677 VSS.n14902 VSS.n14811 0.296
R19678 VSS.n15146 VSS.n15067 0.296
R19679 VSS.n15390 VSS.n15311 0.296
R19680 VSS.n15634 VSS.n15555 0.296
R19681 VSS.n15878 VSS.n15799 0.296
R19682 VSS.n16122 VSS.n16043 0.296
R19683 VSS.n16378 VSS.n16287 0.296
R19684 VSS.n10951 VSS.n10860 0.296
R19685 VSS.n11195 VSS.n11116 0.296
R19686 VSS.n11439 VSS.n11360 0.296
R19687 VSS.n11683 VSS.n11604 0.296
R19688 VSS.n11927 VSS.n11848 0.296
R19689 VSS.n12171 VSS.n12092 0.296
R19690 VSS.n12427 VSS.n12336 0.296
R19691 VSS.n7519 VSS.n7428 0.296
R19692 VSS.n7763 VSS.n7684 0.296
R19693 VSS.n8007 VSS.n7928 0.296
R19694 VSS.n8251 VSS.n8172 0.296
R19695 VSS.n8495 VSS.n8416 0.296
R19696 VSS.n8739 VSS.n8660 0.296
R19697 VSS.n8995 VSS.n8904 0.296
R19698 VSS.n3716 VSS.n3715 0.296
R19699 VSS.n3953 VSS.n3382 0.296
R19700 VSS.n4414 VSS.n4412 0.296
R19701 VSS.n4320 VSS.n4319 0.296
R19702 VSS.n4544 VSS.n3219 0.296
R19703 VSS.n5021 VSS.n4649 0.296
R19704 VSS.n4929 VSS.n4928 0.296
R19705 VSS.n5407 VSS.n1522 0.296
R19706 VSS.n5302 VSS.n1447 0.296
R19707 VSS.n5615 VSS.n1381 0.296
R19708 VSS.n5703 VSS.n589 0.296
R19709 VSS.n883 VSS.n712 0.296
R19710 VSS.n1263 VSS.n1261 0.296
R19711 VSS VSS.n438 0.293
R19712 VSS.n14903 VSS.n14902 0.29
R19713 VSS.n15147 VSS.n15146 0.29
R19714 VSS.n15391 VSS.n15390 0.29
R19715 VSS.n15635 VSS.n15634 0.29
R19716 VSS.n15879 VSS.n15878 0.29
R19717 VSS.n16123 VSS.n16122 0.29
R19718 VSS.n16379 VSS.n16378 0.29
R19719 VSS.n10952 VSS.n10951 0.29
R19720 VSS.n11196 VSS.n11195 0.29
R19721 VSS.n11440 VSS.n11439 0.29
R19722 VSS.n11684 VSS.n11683 0.29
R19723 VSS.n11928 VSS.n11927 0.29
R19724 VSS.n12172 VSS.n12171 0.29
R19725 VSS.n12428 VSS.n12427 0.29
R19726 VSS.n7520 VSS.n7519 0.29
R19727 VSS.n7764 VSS.n7763 0.29
R19728 VSS.n8008 VSS.n8007 0.29
R19729 VSS.n8252 VSS.n8251 0.29
R19730 VSS.n8496 VSS.n8495 0.29
R19731 VSS.n8740 VSS.n8739 0.29
R19732 VSS.n8996 VSS.n8995 0.29
R19733 VSS.n3715 VSS.n3714 0.29
R19734 VSS.n3965 VSS.n3382 0.29
R19735 VSS.n4412 VSS.n4411 0.29
R19736 VSS.n4319 VSS.n4318 0.29
R19737 VSS.n4545 VSS.n4544 0.29
R19738 VSS.n5021 VSS.n5020 0.29
R19739 VSS.n4928 VSS.n4927 0.29
R19740 VSS.n5395 VSS.n1522 0.29
R19741 VSS.n1447 VSS.n1442 0.29
R19742 VSS.n5603 VSS.n1381 0.29
R19743 VSS.n779 VSS.n589 0.29
R19744 VSS.n923 VSS.n712 0.29
R19745 VSS.n1261 VSS.n1260 0.29
R19746 VSS.n16570 VSS.n16527 0.258
R19747 VSS.n12619 VSS.n12576 0.258
R19748 VSS.n9187 VSS.n9144 0.258
R19749 VSS.n1167 VSS.n1166 0.258
R19750 VSS.n5129 VSS.n3096 0.258
R19751 VSS.n18263 VSS.n0 0.256
R19752 VSS.n261 VSS.n260 0.256
R19753 VSS.n18327 VSS.n18326 0.256
R19754 VSS.n243 VSS.n242 0.217
R19755 VSS.n18045 VSS.n18044 0.217
R19756 VSS.n18050 VSS.n18049 0.217
R19757 VSS.n18055 VSS.n18054 0.217
R19758 VSS.n18060 VSS.n18059 0.217
R19759 VSS.n18065 VSS.n18064 0.217
R19760 VSS.n18070 VSS.n18069 0.217
R19761 VSS.n18075 VSS.n18074 0.217
R19762 VSS.n18080 VSS.n18079 0.217
R19763 VSS.n39 VSS.n38 0.217
R19764 VSS.n18261 VSS.n18260 0.217
R19765 VSS.n295 VSS.n294 0.217
R19766 VSS.n17725 VSS.n17724 0.217
R19767 VSS.n17715 VSS.n17714 0.217
R19768 VSS.n17704 VSS.n17703 0.217
R19769 VSS.n17693 VSS.n17692 0.217
R19770 VSS.n17682 VSS.n17681 0.217
R19771 VSS.n17672 VSS.n17671 0.217
R19772 VSS.n17661 VSS.n17660 0.217
R19773 VSS.n17651 VSS.n17650 0.217
R19774 VSS.n18105 VSS.n18104 0.217
R19775 VSS.n18108 VSS.n18107 0.217
R19776 VSS.n17598 VSS.n17597 0.216
R19777 VSS VSS.n14100 0.209
R19778 VSS.n14097 VSS.n14096 0.203
R19779 VSS.t200 VSS.n481 0.201
R19780 VSS.n329 VSS.t180 0.201
R19781 VSS.n17744 VSS.t140 0.201
R19782 VSS.n409 VSS.n359 0.19
R19783 VSS.n410 VSS.n409 0.19
R19784 VSS.n18201 VSS.n18151 0.19
R19785 VSS.n18202 VSS.n18201 0.19
R19786 VSS.n487 VSS.n486 0.178
R19787 VSS.n488 VSS.n487 0.178
R19788 VSS.n489 VSS.n488 0.178
R19789 VSS.n490 VSS.n489 0.178
R19790 VSS.n491 VSS.n490 0.178
R19791 VSS.n474 VSS.n473 0.178
R19792 VSS.n475 VSS.n474 0.178
R19793 VSS.n476 VSS.n475 0.178
R19794 VSS.n477 VSS.n476 0.178
R19795 VSS.n478 VSS.n477 0.178
R19796 VSS.n479 VSS.n478 0.178
R19797 VSS.n480 VSS.n479 0.178
R19798 VSS.n481 VSS.n480 0.178
R19799 VSS.n483 VSS.n482 0.178
R19800 VSS.n484 VSS.n483 0.178
R19801 VSS.n485 VSS.n484 0.178
R19802 VSS.n323 VSS.n322 0.178
R19803 VSS.n324 VSS.n323 0.178
R19804 VSS.n325 VSS.n324 0.178
R19805 VSS.n326 VSS.n325 0.178
R19806 VSS.n327 VSS.n326 0.178
R19807 VSS.n328 VSS.n327 0.178
R19808 VSS.n330 VSS.n329 0.178
R19809 VSS.n17763 VSS.n17762 0.178
R19810 VSS.n17745 VSS.n17744 0.178
R19811 VSS.n17746 VSS.n17745 0.178
R19812 VSS.n17747 VSS.n17746 0.178
R19813 VSS.n17748 VSS.n17747 0.178
R19814 VSS.n17749 VSS.n17748 0.178
R19815 VSS.n17750 VSS.n17749 0.178
R19816 VSS.n17751 VSS.n17750 0.178
R19817 VSS.n17752 VSS.n17751 0.178
R19818 VSS.n17755 VSS.n17754 0.178
R19819 VSS.n17756 VSS.n17755 0.178
R19820 VSS.n17757 VSS.n17756 0.178
R19821 VSS.n17758 VSS.n17757 0.178
R19822 VSS.n17759 VSS.n17758 0.178
R19823 VSS.n17760 VSS.n17759 0.178
R19824 VSS.n17761 VSS.n17760 0.178
R19825 VSS.n10563 VSS.n10562 0.177
R19826 VSS.n18229 VSS.n18228 0.163
R19827 VSS.n331 VSS.n328 0.15
R19828 VSS.n16572 VSS.n16571 0.148
R19829 VSS.n14299 VSS.n14285 0.148
R19830 VSS.n14479 VSS.n14465 0.148
R19831 VSS.n17431 VSS.n17430 0.148
R19832 VSS.n17263 VSS.n17262 0.148
R19833 VSS.n17095 VSS.n17094 0.148
R19834 VSS.n16927 VSS.n16926 0.148
R19835 VSS.n16759 VSS.n16758 0.148
R19836 VSS.n16591 VSS.n16590 0.148
R19837 VSS.n12621 VSS.n12620 0.148
R19838 VSS.n12816 VSS.n12802 0.148
R19839 VSS.n12996 VSS.n12982 0.148
R19840 VSS.n13176 VSS.n13162 0.148
R19841 VSS.n13356 VSS.n13342 0.148
R19842 VSS.n13536 VSS.n13522 0.148
R19843 VSS.n13716 VSS.n13702 0.148
R19844 VSS.n13896 VSS.n13882 0.148
R19845 VSS.n9189 VSS.n9188 0.148
R19846 VSS.n10396 VSS.n10395 0.148
R19847 VSS.n10229 VSS.n10228 0.148
R19848 VSS.n10061 VSS.n10060 0.148
R19849 VSS.n9893 VSS.n9892 0.148
R19850 VSS.n9725 VSS.n9724 0.148
R19851 VSS.n9557 VSS.n9556 0.148
R19852 VSS.n9389 VSS.n9388 0.148
R19853 VSS.n9221 VSS.n9220 0.148
R19854 VSS.n5130 VSS.n3095 0.148
R19855 VSS.n2463 VSS.n2285 0.148
R19856 VSS.n2553 VSS.n2195 0.148
R19857 VSS.n2643 VSS.n2105 0.148
R19858 VSS.n2733 VSS.n2015 0.148
R19859 VSS.n2823 VSS.n1925 0.148
R19860 VSS.n2913 VSS.n1835 0.148
R19861 VSS.n3003 VSS.n1745 0.148
R19862 VSS.n3093 VSS.n1655 0.148
R19863 VSS.n1169 VSS.n1168 0.148
R19864 VSS.n6757 VSS.n6579 0.148
R19865 VSS.n6847 VSS.n6489 0.148
R19866 VSS.n6937 VSS.n6399 0.148
R19867 VSS.n6381 VSS.n5840 0.148
R19868 VSS.n6370 VSS.n6317 0.148
R19869 VSS.n6306 VSS.n6253 0.148
R19870 VSS.n6242 VSS.n6189 0.148
R19871 VSS.n492 VSS.n485 0.148
R19872 VSS.n382 VSS.n381 0.144
R19873 VSS.n389 VSS.n388 0.144
R19874 VSS.n399 VSS.n398 0.144
R19875 VSS.n417 VSS.n416 0.144
R19876 VSS.n424 VSS.n423 0.144
R19877 VSS.n432 VSS.n431 0.144
R19878 VSS.n18174 VSS.n18173 0.144
R19879 VSS.n18181 VSS.n18180 0.144
R19880 VSS.n18191 VSS.n18190 0.144
R19881 VSS.n18210 VSS.n18208 0.144
R19882 VSS.n18217 VSS.n18141 0.144
R19883 VSS.n18219 VSS.n18138 0.144
R19884 VSS.n14313 VSS.n14312 0.142
R19885 VSS.n17597 VSS.n17585 0.142
R19886 VSS.n17429 VSS.n17417 0.142
R19887 VSS.n17261 VSS.n17249 0.142
R19888 VSS.n17093 VSS.n17081 0.142
R19889 VSS.n16925 VSS.n16913 0.142
R19890 VSS.n16757 VSS.n16745 0.142
R19891 VSS.n12830 VSS.n12829 0.142
R19892 VSS.n13010 VSS.n13009 0.142
R19893 VSS.n13190 VSS.n13189 0.142
R19894 VSS.n13370 VSS.n13369 0.142
R19895 VSS.n13550 VSS.n13549 0.142
R19896 VSS.n13730 VSS.n13729 0.142
R19897 VSS.n13910 VSS.n13909 0.142
R19898 VSS.n10382 VSS.n10381 0.142
R19899 VSS.n10214 VSS.n10213 0.142
R19900 VSS.n10046 VSS.n10045 0.142
R19901 VSS.n9878 VSS.n9877 0.142
R19902 VSS.n9710 VSS.n9709 0.142
R19903 VSS.n9542 VSS.n9541 0.142
R19904 VSS.n9374 VSS.n9373 0.142
R19905 VSS.n2464 VSS.n2236 0.142
R19906 VSS.n2554 VSS.n2146 0.142
R19907 VSS.n2644 VSS.n2056 0.142
R19908 VSS.n2734 VSS.n1966 0.142
R19909 VSS.n2824 VSS.n1876 0.142
R19910 VSS.n2914 VSS.n1786 0.142
R19911 VSS.n3004 VSS.n1696 0.142
R19912 VSS.n5133 VSS.n1583 0.142
R19913 VSS.n6758 VSS.n6530 0.142
R19914 VSS.n6848 VSS.n6440 0.142
R19915 VSS.n6380 VSS.n5841 0.142
R19916 VSS.n6316 VSS.n5957 0.142
R19917 VSS.n6252 VSS.n6073 0.142
R19918 VSS.n14063 VSS.n14062 0.132
R19919 VSS.n14661 VSS.n14660 0.13
R19920 VSS.n14675 VSS.n14674 0.13
R19921 VSS.n14689 VSS.n14688 0.13
R19922 VSS.n14703 VSS.n14702 0.13
R19923 VSS.n14717 VSS.n14716 0.13
R19924 VSS.n14738 VSS.n14735 0.13
R19925 VSS.n14736 VSS.n14594 0.13
R19926 VSS.n14753 VSS.n14752 0.13
R19927 VSS.n14767 VSS.n14766 0.13
R19928 VSS.n14781 VSS.n14780 0.13
R19929 VSS.n14795 VSS.n14794 0.13
R19930 VSS.n14917 VSS.n14916 0.13
R19931 VSS.n14931 VSS.n14930 0.13
R19932 VSS.n14945 VSS.n14944 0.13
R19933 VSS.n14959 VSS.n14958 0.13
R19934 VSS.n14973 VSS.n14972 0.13
R19935 VSS.n14994 VSS.n14991 0.13
R19936 VSS.n14992 VSS.n14588 0.13
R19937 VSS.n15009 VSS.n15008 0.13
R19938 VSS.n15023 VSS.n15022 0.13
R19939 VSS.n15037 VSS.n15036 0.13
R19940 VSS.n15051 VSS.n15050 0.13
R19941 VSS.n15161 VSS.n15160 0.13
R19942 VSS.n15175 VSS.n15174 0.13
R19943 VSS.n15189 VSS.n15188 0.13
R19944 VSS.n15203 VSS.n15202 0.13
R19945 VSS.n15217 VSS.n15216 0.13
R19946 VSS.n15238 VSS.n15235 0.13
R19947 VSS.n15236 VSS.n14582 0.13
R19948 VSS.n15253 VSS.n15252 0.13
R19949 VSS.n15267 VSS.n15266 0.13
R19950 VSS.n15281 VSS.n15280 0.13
R19951 VSS.n15295 VSS.n15294 0.13
R19952 VSS.n15405 VSS.n15404 0.13
R19953 VSS.n15419 VSS.n15418 0.13
R19954 VSS.n15433 VSS.n15432 0.13
R19955 VSS.n15447 VSS.n15446 0.13
R19956 VSS.n15461 VSS.n15460 0.13
R19957 VSS.n15482 VSS.n15479 0.13
R19958 VSS.n15480 VSS.n14576 0.13
R19959 VSS.n15497 VSS.n15496 0.13
R19960 VSS.n15511 VSS.n15510 0.13
R19961 VSS.n15525 VSS.n15524 0.13
R19962 VSS.n15539 VSS.n15538 0.13
R19963 VSS.n15649 VSS.n15648 0.13
R19964 VSS.n15663 VSS.n15662 0.13
R19965 VSS.n15677 VSS.n15676 0.13
R19966 VSS.n15691 VSS.n15690 0.13
R19967 VSS.n15705 VSS.n15704 0.13
R19968 VSS.n15726 VSS.n15723 0.13
R19969 VSS.n15724 VSS.n14570 0.13
R19970 VSS.n15741 VSS.n15740 0.13
R19971 VSS.n15755 VSS.n15754 0.13
R19972 VSS.n15769 VSS.n15768 0.13
R19973 VSS.n15783 VSS.n15782 0.13
R19974 VSS.n15893 VSS.n15892 0.13
R19975 VSS.n15907 VSS.n15906 0.13
R19976 VSS.n15921 VSS.n15920 0.13
R19977 VSS.n15935 VSS.n15934 0.13
R19978 VSS.n15949 VSS.n15948 0.13
R19979 VSS.n15970 VSS.n15967 0.13
R19980 VSS.n15968 VSS.n14564 0.13
R19981 VSS.n15985 VSS.n15984 0.13
R19982 VSS.n15999 VSS.n15998 0.13
R19983 VSS.n16013 VSS.n16012 0.13
R19984 VSS.n16027 VSS.n16026 0.13
R19985 VSS.n16137 VSS.n16136 0.13
R19986 VSS.n16151 VSS.n16150 0.13
R19987 VSS.n16165 VSS.n16164 0.13
R19988 VSS.n16179 VSS.n16178 0.13
R19989 VSS.n16193 VSS.n16192 0.13
R19990 VSS.n16214 VSS.n16211 0.13
R19991 VSS.n16212 VSS.n14558 0.13
R19992 VSS.n16229 VSS.n16228 0.13
R19993 VSS.n16243 VSS.n16242 0.13
R19994 VSS.n16257 VSS.n16256 0.13
R19995 VSS.n16271 VSS.n16270 0.13
R19996 VSS.n16393 VSS.n16392 0.13
R19997 VSS.n16407 VSS.n16406 0.13
R19998 VSS.n16421 VSS.n16420 0.13
R19999 VSS.n16435 VSS.n16434 0.13
R20000 VSS.n16449 VSS.n16448 0.13
R20001 VSS.n16470 VSS.n16467 0.13
R20002 VSS.n16468 VSS.n14552 0.13
R20003 VSS.n16485 VSS.n16484 0.13
R20004 VSS.n16499 VSS.n16498 0.13
R20005 VSS.n16513 VSS.n16512 0.13
R20006 VSS.n14145 VSS.n14144 0.13
R20007 VSS.n14157 VSS.n14156 0.13
R20008 VSS.n14169 VSS.n14168 0.13
R20009 VSS.n14181 VSS.n14180 0.13
R20010 VSS.n14193 VSS.n14192 0.13
R20011 VSS.n14205 VSS.n14204 0.13
R20012 VSS.n14217 VSS.n14216 0.13
R20013 VSS.n14229 VSS.n14228 0.13
R20014 VSS.n14325 VSS.n14324 0.13
R20015 VSS.n14337 VSS.n14336 0.13
R20016 VSS.n14349 VSS.n14348 0.13
R20017 VSS.n14361 VSS.n14360 0.13
R20018 VSS.n14373 VSS.n14372 0.13
R20019 VSS.n14385 VSS.n14384 0.13
R20020 VSS.n14397 VSS.n14396 0.13
R20021 VSS.n14409 VSS.n14408 0.13
R20022 VSS.n17527 VSS.n17526 0.13
R20023 VSS.n17515 VSS.n17514 0.13
R20024 VSS.n17503 VSS.n17502 0.13
R20025 VSS.n17491 VSS.n17490 0.13
R20026 VSS.n17479 VSS.n17478 0.13
R20027 VSS.n17467 VSS.n17466 0.13
R20028 VSS.n17455 VSS.n17454 0.13
R20029 VSS.n17443 VSS.n17442 0.13
R20030 VSS.n17359 VSS.n17358 0.13
R20031 VSS.n17347 VSS.n17346 0.13
R20032 VSS.n17335 VSS.n17334 0.13
R20033 VSS.n17323 VSS.n17322 0.13
R20034 VSS.n17311 VSS.n17310 0.13
R20035 VSS.n17299 VSS.n17298 0.13
R20036 VSS.n17287 VSS.n17286 0.13
R20037 VSS.n17275 VSS.n17274 0.13
R20038 VSS.n17191 VSS.n17190 0.13
R20039 VSS.n17179 VSS.n17178 0.13
R20040 VSS.n17167 VSS.n17166 0.13
R20041 VSS.n17155 VSS.n17154 0.13
R20042 VSS.n17143 VSS.n17142 0.13
R20043 VSS.n17131 VSS.n17130 0.13
R20044 VSS.n17119 VSS.n17118 0.13
R20045 VSS.n17107 VSS.n17106 0.13
R20046 VSS.n17023 VSS.n17022 0.13
R20047 VSS.n17011 VSS.n17010 0.13
R20048 VSS.n16999 VSS.n16998 0.13
R20049 VSS.n16987 VSS.n16986 0.13
R20050 VSS.n16975 VSS.n16974 0.13
R20051 VSS.n16963 VSS.n16962 0.13
R20052 VSS.n16951 VSS.n16950 0.13
R20053 VSS.n16939 VSS.n16938 0.13
R20054 VSS.n16855 VSS.n16854 0.13
R20055 VSS.n16843 VSS.n16842 0.13
R20056 VSS.n16831 VSS.n16830 0.13
R20057 VSS.n16819 VSS.n16818 0.13
R20058 VSS.n16807 VSS.n16806 0.13
R20059 VSS.n16795 VSS.n16794 0.13
R20060 VSS.n16783 VSS.n16782 0.13
R20061 VSS.n16771 VSS.n16770 0.13
R20062 VSS.n16687 VSS.n16686 0.13
R20063 VSS.n16675 VSS.n16674 0.13
R20064 VSS.n16663 VSS.n16662 0.13
R20065 VSS.n16651 VSS.n16650 0.13
R20066 VSS.n16639 VSS.n16638 0.13
R20067 VSS.n16627 VSS.n16626 0.13
R20068 VSS.n16615 VSS.n16614 0.13
R20069 VSS.n16603 VSS.n16602 0.13
R20070 VSS.n10710 VSS.n10709 0.13
R20071 VSS.n10724 VSS.n10723 0.13
R20072 VSS.n10738 VSS.n10737 0.13
R20073 VSS.n10752 VSS.n10751 0.13
R20074 VSS.n10766 VSS.n10765 0.13
R20075 VSS.n10787 VSS.n10784 0.13
R20076 VSS.n10785 VSS.n10643 0.13
R20077 VSS.n10802 VSS.n10801 0.13
R20078 VSS.n10816 VSS.n10815 0.13
R20079 VSS.n10830 VSS.n10829 0.13
R20080 VSS.n10844 VSS.n10843 0.13
R20081 VSS.n10966 VSS.n10965 0.13
R20082 VSS.n10980 VSS.n10979 0.13
R20083 VSS.n10994 VSS.n10993 0.13
R20084 VSS.n11008 VSS.n11007 0.13
R20085 VSS.n11022 VSS.n11021 0.13
R20086 VSS.n11043 VSS.n11040 0.13
R20087 VSS.n11041 VSS.n10637 0.13
R20088 VSS.n11058 VSS.n11057 0.13
R20089 VSS.n11072 VSS.n11071 0.13
R20090 VSS.n11086 VSS.n11085 0.13
R20091 VSS.n11100 VSS.n11099 0.13
R20092 VSS.n11210 VSS.n11209 0.13
R20093 VSS.n11224 VSS.n11223 0.13
R20094 VSS.n11238 VSS.n11237 0.13
R20095 VSS.n11252 VSS.n11251 0.13
R20096 VSS.n11266 VSS.n11265 0.13
R20097 VSS.n11287 VSS.n11284 0.13
R20098 VSS.n11285 VSS.n10631 0.13
R20099 VSS.n11302 VSS.n11301 0.13
R20100 VSS.n11316 VSS.n11315 0.13
R20101 VSS.n11330 VSS.n11329 0.13
R20102 VSS.n11344 VSS.n11343 0.13
R20103 VSS.n11454 VSS.n11453 0.13
R20104 VSS.n11468 VSS.n11467 0.13
R20105 VSS.n11482 VSS.n11481 0.13
R20106 VSS.n11496 VSS.n11495 0.13
R20107 VSS.n11510 VSS.n11509 0.13
R20108 VSS.n11531 VSS.n11528 0.13
R20109 VSS.n11529 VSS.n10625 0.13
R20110 VSS.n11546 VSS.n11545 0.13
R20111 VSS.n11560 VSS.n11559 0.13
R20112 VSS.n11574 VSS.n11573 0.13
R20113 VSS.n11588 VSS.n11587 0.13
R20114 VSS.n11698 VSS.n11697 0.13
R20115 VSS.n11712 VSS.n11711 0.13
R20116 VSS.n11726 VSS.n11725 0.13
R20117 VSS.n11740 VSS.n11739 0.13
R20118 VSS.n11754 VSS.n11753 0.13
R20119 VSS.n11775 VSS.n11772 0.13
R20120 VSS.n11773 VSS.n10619 0.13
R20121 VSS.n11790 VSS.n11789 0.13
R20122 VSS.n11804 VSS.n11803 0.13
R20123 VSS.n11818 VSS.n11817 0.13
R20124 VSS.n11832 VSS.n11831 0.13
R20125 VSS.n11942 VSS.n11941 0.13
R20126 VSS.n11956 VSS.n11955 0.13
R20127 VSS.n11970 VSS.n11969 0.13
R20128 VSS.n11984 VSS.n11983 0.13
R20129 VSS.n11998 VSS.n11997 0.13
R20130 VSS.n12019 VSS.n12016 0.13
R20131 VSS.n12017 VSS.n10613 0.13
R20132 VSS.n12034 VSS.n12033 0.13
R20133 VSS.n12048 VSS.n12047 0.13
R20134 VSS.n12062 VSS.n12061 0.13
R20135 VSS.n12076 VSS.n12075 0.13
R20136 VSS.n12186 VSS.n12185 0.13
R20137 VSS.n12200 VSS.n12199 0.13
R20138 VSS.n12214 VSS.n12213 0.13
R20139 VSS.n12228 VSS.n12227 0.13
R20140 VSS.n12242 VSS.n12241 0.13
R20141 VSS.n12263 VSS.n12260 0.13
R20142 VSS.n12261 VSS.n10607 0.13
R20143 VSS.n12278 VSS.n12277 0.13
R20144 VSS.n12292 VSS.n12291 0.13
R20145 VSS.n12306 VSS.n12305 0.13
R20146 VSS.n12320 VSS.n12319 0.13
R20147 VSS.n12442 VSS.n12441 0.13
R20148 VSS.n12456 VSS.n12455 0.13
R20149 VSS.n12470 VSS.n12469 0.13
R20150 VSS.n12484 VSS.n12483 0.13
R20151 VSS.n12498 VSS.n12497 0.13
R20152 VSS.n12519 VSS.n12516 0.13
R20153 VSS.n12517 VSS.n10601 0.13
R20154 VSS.n12534 VSS.n12533 0.13
R20155 VSS.n12548 VSS.n12547 0.13
R20156 VSS.n12562 VSS.n12561 0.13
R20157 VSS.n12662 VSS.n12661 0.13
R20158 VSS.n12674 VSS.n12673 0.13
R20159 VSS.n12686 VSS.n12685 0.13
R20160 VSS.n12698 VSS.n12697 0.13
R20161 VSS.n12710 VSS.n12709 0.13
R20162 VSS.n12722 VSS.n12721 0.13
R20163 VSS.n12734 VSS.n12733 0.13
R20164 VSS.n12746 VSS.n12745 0.13
R20165 VSS.n12842 VSS.n12841 0.13
R20166 VSS.n12854 VSS.n12853 0.13
R20167 VSS.n12866 VSS.n12865 0.13
R20168 VSS.n12878 VSS.n12877 0.13
R20169 VSS.n12890 VSS.n12889 0.13
R20170 VSS.n12902 VSS.n12901 0.13
R20171 VSS.n12914 VSS.n12913 0.13
R20172 VSS.n12926 VSS.n12925 0.13
R20173 VSS.n13022 VSS.n13021 0.13
R20174 VSS.n13034 VSS.n13033 0.13
R20175 VSS.n13046 VSS.n13045 0.13
R20176 VSS.n13058 VSS.n13057 0.13
R20177 VSS.n13070 VSS.n13069 0.13
R20178 VSS.n13082 VSS.n13081 0.13
R20179 VSS.n13094 VSS.n13093 0.13
R20180 VSS.n13106 VSS.n13105 0.13
R20181 VSS.n13202 VSS.n13201 0.13
R20182 VSS.n13214 VSS.n13213 0.13
R20183 VSS.n13226 VSS.n13225 0.13
R20184 VSS.n13238 VSS.n13237 0.13
R20185 VSS.n13250 VSS.n13249 0.13
R20186 VSS.n13262 VSS.n13261 0.13
R20187 VSS.n13274 VSS.n13273 0.13
R20188 VSS.n13286 VSS.n13285 0.13
R20189 VSS.n13382 VSS.n13381 0.13
R20190 VSS.n13394 VSS.n13393 0.13
R20191 VSS.n13406 VSS.n13405 0.13
R20192 VSS.n13418 VSS.n13417 0.13
R20193 VSS.n13430 VSS.n13429 0.13
R20194 VSS.n13442 VSS.n13441 0.13
R20195 VSS.n13454 VSS.n13453 0.13
R20196 VSS.n13466 VSS.n13465 0.13
R20197 VSS.n13562 VSS.n13561 0.13
R20198 VSS.n13574 VSS.n13573 0.13
R20199 VSS.n13586 VSS.n13585 0.13
R20200 VSS.n13598 VSS.n13597 0.13
R20201 VSS.n13610 VSS.n13609 0.13
R20202 VSS.n13622 VSS.n13621 0.13
R20203 VSS.n13634 VSS.n13633 0.13
R20204 VSS.n13646 VSS.n13645 0.13
R20205 VSS.n13742 VSS.n13741 0.13
R20206 VSS.n13754 VSS.n13753 0.13
R20207 VSS.n13766 VSS.n13765 0.13
R20208 VSS.n13778 VSS.n13777 0.13
R20209 VSS.n13790 VSS.n13789 0.13
R20210 VSS.n13802 VSS.n13801 0.13
R20211 VSS.n13814 VSS.n13813 0.13
R20212 VSS.n13826 VSS.n13825 0.13
R20213 VSS.n13922 VSS.n13921 0.13
R20214 VSS.n13934 VSS.n13933 0.13
R20215 VSS.n13946 VSS.n13945 0.13
R20216 VSS.n13958 VSS.n13957 0.13
R20217 VSS.n13970 VSS.n13969 0.13
R20218 VSS.n13982 VSS.n13981 0.13
R20219 VSS.n13994 VSS.n13993 0.13
R20220 VSS.n14006 VSS.n14005 0.13
R20221 VSS.n7278 VSS.n7277 0.13
R20222 VSS.n7292 VSS.n7291 0.13
R20223 VSS.n7306 VSS.n7305 0.13
R20224 VSS.n7320 VSS.n7319 0.13
R20225 VSS.n7334 VSS.n7333 0.13
R20226 VSS.n7355 VSS.n7352 0.13
R20227 VSS.n7353 VSS.n7211 0.13
R20228 VSS.n7370 VSS.n7369 0.13
R20229 VSS.n7384 VSS.n7383 0.13
R20230 VSS.n7398 VSS.n7397 0.13
R20231 VSS.n7412 VSS.n7411 0.13
R20232 VSS.n7534 VSS.n7533 0.13
R20233 VSS.n7548 VSS.n7547 0.13
R20234 VSS.n7562 VSS.n7561 0.13
R20235 VSS.n7576 VSS.n7575 0.13
R20236 VSS.n7590 VSS.n7589 0.13
R20237 VSS.n7611 VSS.n7608 0.13
R20238 VSS.n7609 VSS.n7205 0.13
R20239 VSS.n7626 VSS.n7625 0.13
R20240 VSS.n7640 VSS.n7639 0.13
R20241 VSS.n7654 VSS.n7653 0.13
R20242 VSS.n7668 VSS.n7667 0.13
R20243 VSS.n7778 VSS.n7777 0.13
R20244 VSS.n7792 VSS.n7791 0.13
R20245 VSS.n7806 VSS.n7805 0.13
R20246 VSS.n7820 VSS.n7819 0.13
R20247 VSS.n7834 VSS.n7833 0.13
R20248 VSS.n7855 VSS.n7852 0.13
R20249 VSS.n7853 VSS.n7199 0.13
R20250 VSS.n7870 VSS.n7869 0.13
R20251 VSS.n7884 VSS.n7883 0.13
R20252 VSS.n7898 VSS.n7897 0.13
R20253 VSS.n7912 VSS.n7911 0.13
R20254 VSS.n8022 VSS.n8021 0.13
R20255 VSS.n8036 VSS.n8035 0.13
R20256 VSS.n8050 VSS.n8049 0.13
R20257 VSS.n8064 VSS.n8063 0.13
R20258 VSS.n8078 VSS.n8077 0.13
R20259 VSS.n8099 VSS.n8096 0.13
R20260 VSS.n8097 VSS.n7193 0.13
R20261 VSS.n8114 VSS.n8113 0.13
R20262 VSS.n8128 VSS.n8127 0.13
R20263 VSS.n8142 VSS.n8141 0.13
R20264 VSS.n8156 VSS.n8155 0.13
R20265 VSS.n8266 VSS.n8265 0.13
R20266 VSS.n8280 VSS.n8279 0.13
R20267 VSS.n8294 VSS.n8293 0.13
R20268 VSS.n8308 VSS.n8307 0.13
R20269 VSS.n8322 VSS.n8321 0.13
R20270 VSS.n8343 VSS.n8340 0.13
R20271 VSS.n8341 VSS.n7187 0.13
R20272 VSS.n8358 VSS.n8357 0.13
R20273 VSS.n8372 VSS.n8371 0.13
R20274 VSS.n8386 VSS.n8385 0.13
R20275 VSS.n8400 VSS.n8399 0.13
R20276 VSS.n8510 VSS.n8509 0.13
R20277 VSS.n8524 VSS.n8523 0.13
R20278 VSS.n8538 VSS.n8537 0.13
R20279 VSS.n8552 VSS.n8551 0.13
R20280 VSS.n8566 VSS.n8565 0.13
R20281 VSS.n8587 VSS.n8584 0.13
R20282 VSS.n8585 VSS.n7181 0.13
R20283 VSS.n8602 VSS.n8601 0.13
R20284 VSS.n8616 VSS.n8615 0.13
R20285 VSS.n8630 VSS.n8629 0.13
R20286 VSS.n8644 VSS.n8643 0.13
R20287 VSS.n8754 VSS.n8753 0.13
R20288 VSS.n8768 VSS.n8767 0.13
R20289 VSS.n8782 VSS.n8781 0.13
R20290 VSS.n8796 VSS.n8795 0.13
R20291 VSS.n8810 VSS.n8809 0.13
R20292 VSS.n8831 VSS.n8828 0.13
R20293 VSS.n8829 VSS.n7175 0.13
R20294 VSS.n8846 VSS.n8845 0.13
R20295 VSS.n8860 VSS.n8859 0.13
R20296 VSS.n8874 VSS.n8873 0.13
R20297 VSS.n8888 VSS.n8887 0.13
R20298 VSS.n9010 VSS.n9009 0.13
R20299 VSS.n9024 VSS.n9023 0.13
R20300 VSS.n9038 VSS.n9037 0.13
R20301 VSS.n9052 VSS.n9051 0.13
R20302 VSS.n9066 VSS.n9065 0.13
R20303 VSS.n9087 VSS.n9084 0.13
R20304 VSS.n9085 VSS.n7169 0.13
R20305 VSS.n9102 VSS.n9101 0.13
R20306 VSS.n9116 VSS.n9115 0.13
R20307 VSS.n9130 VSS.n9129 0.13
R20308 VSS.n10492 VSS.n10491 0.13
R20309 VSS.n10480 VSS.n10479 0.13
R20310 VSS.n10468 VSS.n10467 0.13
R20311 VSS.n10456 VSS.n10455 0.13
R20312 VSS.n10444 VSS.n10443 0.13
R20313 VSS.n10432 VSS.n10431 0.13
R20314 VSS.n10420 VSS.n10419 0.13
R20315 VSS.n10408 VSS.n10407 0.13
R20316 VSS.n10325 VSS.n10324 0.13
R20317 VSS.n10313 VSS.n10312 0.13
R20318 VSS.n10301 VSS.n10300 0.13
R20319 VSS.n10289 VSS.n10288 0.13
R20320 VSS.n10277 VSS.n10276 0.13
R20321 VSS.n10265 VSS.n10264 0.13
R20322 VSS.n10253 VSS.n10252 0.13
R20323 VSS.n10241 VSS.n10240 0.13
R20324 VSS.n10157 VSS.n10156 0.13
R20325 VSS.n10145 VSS.n10144 0.13
R20326 VSS.n10133 VSS.n10132 0.13
R20327 VSS.n10121 VSS.n10120 0.13
R20328 VSS.n10109 VSS.n10108 0.13
R20329 VSS.n10097 VSS.n10096 0.13
R20330 VSS.n10085 VSS.n10084 0.13
R20331 VSS.n10073 VSS.n10072 0.13
R20332 VSS.n9989 VSS.n9988 0.13
R20333 VSS.n9977 VSS.n9976 0.13
R20334 VSS.n9965 VSS.n9964 0.13
R20335 VSS.n9953 VSS.n9952 0.13
R20336 VSS.n9941 VSS.n9940 0.13
R20337 VSS.n9929 VSS.n9928 0.13
R20338 VSS.n9917 VSS.n9916 0.13
R20339 VSS.n9905 VSS.n9904 0.13
R20340 VSS.n9821 VSS.n9820 0.13
R20341 VSS.n9809 VSS.n9808 0.13
R20342 VSS.n9797 VSS.n9796 0.13
R20343 VSS.n9785 VSS.n9784 0.13
R20344 VSS.n9773 VSS.n9772 0.13
R20345 VSS.n9761 VSS.n9760 0.13
R20346 VSS.n9749 VSS.n9748 0.13
R20347 VSS.n9737 VSS.n9736 0.13
R20348 VSS.n9653 VSS.n9652 0.13
R20349 VSS.n9641 VSS.n9640 0.13
R20350 VSS.n9629 VSS.n9628 0.13
R20351 VSS.n9617 VSS.n9616 0.13
R20352 VSS.n9605 VSS.n9604 0.13
R20353 VSS.n9593 VSS.n9592 0.13
R20354 VSS.n9581 VSS.n9580 0.13
R20355 VSS.n9569 VSS.n9568 0.13
R20356 VSS.n9485 VSS.n9484 0.13
R20357 VSS.n9473 VSS.n9472 0.13
R20358 VSS.n9461 VSS.n9460 0.13
R20359 VSS.n9449 VSS.n9448 0.13
R20360 VSS.n9437 VSS.n9436 0.13
R20361 VSS.n9425 VSS.n9424 0.13
R20362 VSS.n9413 VSS.n9412 0.13
R20363 VSS.n9401 VSS.n9400 0.13
R20364 VSS.n9317 VSS.n9316 0.13
R20365 VSS.n9305 VSS.n9304 0.13
R20366 VSS.n9293 VSS.n9292 0.13
R20367 VSS.n9281 VSS.n9280 0.13
R20368 VSS.n9269 VSS.n9268 0.13
R20369 VSS.n9257 VSS.n9256 0.13
R20370 VSS.n9245 VSS.n9244 0.13
R20371 VSS.n9233 VSS.n9232 0.13
R20372 VSS.n3798 VSS.n3461 0.13
R20373 VSS.n3796 VSS.n3462 0.13
R20374 VSS.n3785 VSS.n3784 0.13
R20375 VSS.n3775 VSS.n3480 0.13
R20376 VSS.n3773 VSS.n3481 0.13
R20377 VSS.n3762 VSS.n3761 0.13
R20378 VSS.n3752 VSS.n3499 0.13
R20379 VSS.n3750 VSS.n3500 0.13
R20380 VSS.n3739 VSS.n3738 0.13
R20381 VSS.n3729 VSS.n3518 0.13
R20382 VSS.n3727 VSS.n3519 0.13
R20383 VSS.n3705 VSS.n3573 0.13
R20384 VSS.n3703 VSS.n3574 0.13
R20385 VSS.n3692 VSS.n3691 0.13
R20386 VSS.n3682 VSS.n3592 0.13
R20387 VSS.n3680 VSS.n3593 0.13
R20388 VSS.n3669 VSS.n3668 0.13
R20389 VSS.n3659 VSS.n3611 0.13
R20390 VSS.n3657 VSS.n3612 0.13
R20391 VSS.n3646 VSS.n3645 0.13
R20392 VSS.n3636 VSS.n3634 0.13
R20393 VSS.n3955 VSS.n3391 0.13
R20394 VSS.n3967 VSS.n3377 0.13
R20395 VSS.n3979 VSS.n3978 0.13
R20396 VSS.n3991 VSS.n3989 0.13
R20397 VSS.n4000 VSS.n3361 0.13
R20398 VSS.n4002 VSS.n3356 0.13
R20399 VSS.n4014 VSS.n4013 0.13
R20400 VSS.n4026 VSS.n4024 0.13
R20401 VSS.n4035 VSS.n3340 0.13
R20402 VSS.n4037 VSS.n3335 0.13
R20403 VSS.n4049 VSS.n4048 0.13
R20404 VSS.n4416 VSS.n4059 0.13
R20405 VSS.n4402 VSS.n4073 0.13
R20406 VSS.n4400 VSS.n4074 0.13
R20407 VSS.n4389 VSS.n4388 0.13
R20408 VSS.n4379 VSS.n4092 0.13
R20409 VSS.n4377 VSS.n4093 0.13
R20410 VSS.n4366 VSS.n4365 0.13
R20411 VSS.n4356 VSS.n4111 0.13
R20412 VSS.n4354 VSS.n4112 0.13
R20413 VSS.n4343 VSS.n4342 0.13
R20414 VSS.n4333 VSS.n4130 0.13
R20415 VSS.n4331 VSS.n4131 0.13
R20416 VSS.n4309 VSS.n4185 0.13
R20417 VSS.n4307 VSS.n4186 0.13
R20418 VSS.n4296 VSS.n4295 0.13
R20419 VSS.n4286 VSS.n4204 0.13
R20420 VSS.n4284 VSS.n4205 0.13
R20421 VSS.n4273 VSS.n4272 0.13
R20422 VSS.n4263 VSS.n4223 0.13
R20423 VSS.n4261 VSS.n4224 0.13
R20424 VSS.n4250 VSS.n4249 0.13
R20425 VSS.n4240 VSS.n4239 0.13
R20426 VSS.n4539 VSS.n4538 0.13
R20427 VSS.n4557 VSS.n4555 0.13
R20428 VSS.n4566 VSS.n3205 0.13
R20429 VSS.n4568 VSS.n3200 0.13
R20430 VSS.n4580 VSS.n4579 0.13
R20431 VSS.n4592 VSS.n4590 0.13
R20432 VSS.n4601 VSS.n3184 0.13
R20433 VSS.n4603 VSS.n3179 0.13
R20434 VSS.n4615 VSS.n4614 0.13
R20435 VSS.n4627 VSS.n4625 0.13
R20436 VSS.n4636 VSS.n3163 0.13
R20437 VSS.n4638 VSS.n3157 0.13
R20438 VSS.n5011 VSS.n4663 0.13
R20439 VSS.n5009 VSS.n4664 0.13
R20440 VSS.n4998 VSS.n4997 0.13
R20441 VSS.n4988 VSS.n4682 0.13
R20442 VSS.n4986 VSS.n4683 0.13
R20443 VSS.n4975 VSS.n4974 0.13
R20444 VSS.n4965 VSS.n4701 0.13
R20445 VSS.n4963 VSS.n4702 0.13
R20446 VSS.n4952 VSS.n4951 0.13
R20447 VSS.n4942 VSS.n4720 0.13
R20448 VSS.n4940 VSS.n4721 0.13
R20449 VSS.n4918 VSS.n4775 0.13
R20450 VSS.n4916 VSS.n4776 0.13
R20451 VSS.n4905 VSS.n4904 0.13
R20452 VSS.n4895 VSS.n4794 0.13
R20453 VSS.n4893 VSS.n4795 0.13
R20454 VSS.n4882 VSS.n4881 0.13
R20455 VSS.n4872 VSS.n4813 0.13
R20456 VSS.n4870 VSS.n4814 0.13
R20457 VSS.n4859 VSS.n4858 0.13
R20458 VSS.n4849 VSS.n4832 0.13
R20459 VSS.n4847 VSS.n4833 0.13
R20460 VSS.n2451 VSS.n2382 0.13
R20461 VSS.n2449 VSS.n2383 0.13
R20462 VSS.n2440 VSS.n2439 0.13
R20463 VSS.n2434 VSS.n2433 0.13
R20464 VSS.n2428 VSS.n2427 0.13
R20465 VSS.n2422 VSS.n2421 0.13
R20466 VSS.n2417 VSS.n2416 0.13
R20467 VSS.n2411 VSS.n2410 0.13
R20468 VSS.n2541 VSS.n2472 0.13
R20469 VSS.n2539 VSS.n2473 0.13
R20470 VSS.n2530 VSS.n2529 0.13
R20471 VSS.n2524 VSS.n2523 0.13
R20472 VSS.n2518 VSS.n2517 0.13
R20473 VSS.n2512 VSS.n2511 0.13
R20474 VSS.n2507 VSS.n2506 0.13
R20475 VSS.n2501 VSS.n2500 0.13
R20476 VSS.n2631 VSS.n2562 0.13
R20477 VSS.n2629 VSS.n2563 0.13
R20478 VSS.n2620 VSS.n2619 0.13
R20479 VSS.n2614 VSS.n2613 0.13
R20480 VSS.n2608 VSS.n2607 0.13
R20481 VSS.n2602 VSS.n2601 0.13
R20482 VSS.n2597 VSS.n2596 0.13
R20483 VSS.n2591 VSS.n2590 0.13
R20484 VSS.n2721 VSS.n2652 0.13
R20485 VSS.n2719 VSS.n2653 0.13
R20486 VSS.n2710 VSS.n2709 0.13
R20487 VSS.n2704 VSS.n2703 0.13
R20488 VSS.n2698 VSS.n2697 0.13
R20489 VSS.n2692 VSS.n2691 0.13
R20490 VSS.n2687 VSS.n2686 0.13
R20491 VSS.n2681 VSS.n2680 0.13
R20492 VSS.n2811 VSS.n2742 0.13
R20493 VSS.n2809 VSS.n2743 0.13
R20494 VSS.n2800 VSS.n2799 0.13
R20495 VSS.n2794 VSS.n2793 0.13
R20496 VSS.n2788 VSS.n2787 0.13
R20497 VSS.n2782 VSS.n2781 0.13
R20498 VSS.n2777 VSS.n2776 0.13
R20499 VSS.n2771 VSS.n2770 0.13
R20500 VSS.n2901 VSS.n2832 0.13
R20501 VSS.n2899 VSS.n2833 0.13
R20502 VSS.n2890 VSS.n2889 0.13
R20503 VSS.n2884 VSS.n2883 0.13
R20504 VSS.n2878 VSS.n2877 0.13
R20505 VSS.n2872 VSS.n2871 0.13
R20506 VSS.n2867 VSS.n2866 0.13
R20507 VSS.n2861 VSS.n2860 0.13
R20508 VSS.n2991 VSS.n2922 0.13
R20509 VSS.n2989 VSS.n2923 0.13
R20510 VSS.n2980 VSS.n2979 0.13
R20511 VSS.n2974 VSS.n2973 0.13
R20512 VSS.n2968 VSS.n2967 0.13
R20513 VSS.n2962 VSS.n2961 0.13
R20514 VSS.n2957 VSS.n2956 0.13
R20515 VSS.n2951 VSS.n2950 0.13
R20516 VSS.n3081 VSS.n3012 0.13
R20517 VSS.n3079 VSS.n3013 0.13
R20518 VSS.n3070 VSS.n3069 0.13
R20519 VSS.n3064 VSS.n3063 0.13
R20520 VSS.n3058 VSS.n3057 0.13
R20521 VSS.n3052 VSS.n3051 0.13
R20522 VSS.n3047 VSS.n3046 0.13
R20523 VSS.n3041 VSS.n3040 0.13
R20524 VSS.n5145 VSS.n5144 0.13
R20525 VSS.n5157 VSS.n5155 0.13
R20526 VSS.n5166 VSS.n1567 0.13
R20527 VSS.n5168 VSS.n1562 0.13
R20528 VSS.n5180 VSS.n5179 0.13
R20529 VSS.n5192 VSS.n5190 0.13
R20530 VSS.n5201 VSS.n1546 0.13
R20531 VSS.n5203 VSS.n1541 0.13
R20532 VSS.n5215 VSS.n5214 0.13
R20533 VSS.n5227 VSS.n5226 0.13
R20534 VSS.n5405 VSS.n1524 0.13
R20535 VSS.n5393 VSS.n5238 0.13
R20536 VSS.n5382 VSS.n5381 0.13
R20537 VSS.n5372 VSS.n5257 0.13
R20538 VSS.n5370 VSS.n5258 0.13
R20539 VSS.n5359 VSS.n5358 0.13
R20540 VSS.n5349 VSS.n5276 0.13
R20541 VSS.n5347 VSS.n5277 0.13
R20542 VSS.n5336 VSS.n5335 0.13
R20543 VSS.n5326 VSS.n5295 0.13
R20544 VSS.n5324 VSS.n5296 0.13
R20545 VSS.n5313 VSS.n5312 0.13
R20546 VSS.n5504 VSS.n5503 0.13
R20547 VSS.n5516 VSS.n5514 0.13
R20548 VSS.n5525 VSS.n1426 0.13
R20549 VSS.n5527 VSS.n1421 0.13
R20550 VSS.n5539 VSS.n5538 0.13
R20551 VSS.n5551 VSS.n5549 0.13
R20552 VSS.n5560 VSS.n1405 0.13
R20553 VSS.n5562 VSS.n1400 0.13
R20554 VSS.n5574 VSS.n5573 0.13
R20555 VSS.n5586 VSS.n5585 0.13
R20556 VSS.n5613 VSS.n1383 0.13
R20557 VSS.n5774 VSS.n531 0.13
R20558 VSS.n5772 VSS.n532 0.13
R20559 VSS.n5761 VSS.n5760 0.13
R20560 VSS.n5751 VSS.n550 0.13
R20561 VSS.n5749 VSS.n551 0.13
R20562 VSS.n5738 VSS.n5737 0.13
R20563 VSS.n5728 VSS.n569 0.13
R20564 VSS.n5726 VSS.n570 0.13
R20565 VSS.n5715 VSS.n5714 0.13
R20566 VSS.n5705 VSS.n588 0.13
R20567 VSS.n790 VSS.n789 0.13
R20568 VSS.n802 VSS.n800 0.13
R20569 VSS.n811 VSS.n763 0.13
R20570 VSS.n813 VSS.n758 0.13
R20571 VSS.n825 VSS.n824 0.13
R20572 VSS.n837 VSS.n835 0.13
R20573 VSS.n846 VSS.n742 0.13
R20574 VSS.n848 VSS.n737 0.13
R20575 VSS.n860 VSS.n859 0.13
R20576 VSS.n872 VSS.n870 0.13
R20577 VSS.n881 VSS.n720 0.13
R20578 VSS.n925 VSS.n707 0.13
R20579 VSS.n937 VSS.n936 0.13
R20580 VSS.n949 VSS.n947 0.13
R20581 VSS.n958 VSS.n691 0.13
R20582 VSS.n960 VSS.n686 0.13
R20583 VSS.n972 VSS.n971 0.13
R20584 VSS.n984 VSS.n982 0.13
R20585 VSS.n993 VSS.n670 0.13
R20586 VSS.n995 VSS.n665 0.13
R20587 VSS.n1007 VSS.n1006 0.13
R20588 VSS.n1265 VSS.n1017 0.13
R20589 VSS.n1251 VSS.n1031 0.13
R20590 VSS.n1249 VSS.n1032 0.13
R20591 VSS.n1238 VSS.n1237 0.13
R20592 VSS.n1228 VSS.n1050 0.13
R20593 VSS.n1226 VSS.n1051 0.13
R20594 VSS.n1215 VSS.n1214 0.13
R20595 VSS.n1205 VSS.n1069 0.13
R20596 VSS.n1203 VSS.n1070 0.13
R20597 VSS.n1192 VSS.n1191 0.13
R20598 VSS.n1182 VSS.n1088 0.13
R20599 VSS.n1180 VSS.n1089 0.13
R20600 VSS.n6744 VSS.n6676 0.13
R20601 VSS.n6742 VSS.n6677 0.13
R20602 VSS.n6733 VSS.n6732 0.13
R20603 VSS.n6727 VSS.n6726 0.13
R20604 VSS.n6721 VSS.n6720 0.13
R20605 VSS.n6715 VSS.n6714 0.13
R20606 VSS.n6709 VSS.n6708 0.13
R20607 VSS.n6704 VSS.n6703 0.13
R20608 VSS.n6834 VSS.n6766 0.13
R20609 VSS.n6832 VSS.n6767 0.13
R20610 VSS.n6823 VSS.n6822 0.13
R20611 VSS.n6817 VSS.n6816 0.13
R20612 VSS.n6811 VSS.n6810 0.13
R20613 VSS.n6805 VSS.n6804 0.13
R20614 VSS.n6799 VSS.n6798 0.13
R20615 VSS.n6794 VSS.n6793 0.13
R20616 VSS.n6924 VSS.n6856 0.13
R20617 VSS.n6922 VSS.n6857 0.13
R20618 VSS.n6913 VSS.n6912 0.13
R20619 VSS.n6907 VSS.n6906 0.13
R20620 VSS.n6901 VSS.n6900 0.13
R20621 VSS.n6895 VSS.n6894 0.13
R20622 VSS.n6889 VSS.n6888 0.13
R20623 VSS.n6884 VSS.n6883 0.13
R20624 VSS.n5794 VSS.n5793 0.13
R20625 VSS.n5800 VSS.n5799 0.13
R20626 VSS.n5806 VSS.n5805 0.13
R20627 VSS.n5812 VSS.n5811 0.13
R20628 VSS.n5817 VSS.n5816 0.13
R20629 VSS.n5824 VSS.n5823 0.13
R20630 VSS.n5830 VSS.n5829 0.13
R20631 VSS.n5836 VSS.n5835 0.13
R20632 VSS.n5901 VSS.n5900 0.13
R20633 VSS.n5909 VSS.n5908 0.13
R20634 VSS.n5917 VSS.n5916 0.13
R20635 VSS.n5925 VSS.n5924 0.13
R20636 VSS.n5933 VSS.n5932 0.13
R20637 VSS.n5941 VSS.n5940 0.13
R20638 VSS.n5949 VSS.n5948 0.13
R20639 VSS.n6372 VSS.n5956 0.13
R20640 VSS.n6017 VSS.n6016 0.13
R20641 VSS.n6025 VSS.n6024 0.13
R20642 VSS.n6033 VSS.n6032 0.13
R20643 VSS.n6041 VSS.n6040 0.13
R20644 VSS.n6049 VSS.n6048 0.13
R20645 VSS.n6057 VSS.n6056 0.13
R20646 VSS.n6065 VSS.n6064 0.13
R20647 VSS.n6308 VSS.n6072 0.13
R20648 VSS.n6133 VSS.n6132 0.13
R20649 VSS.n6141 VSS.n6140 0.13
R20650 VSS.n6149 VSS.n6148 0.13
R20651 VSS.n6157 VSS.n6156 0.13
R20652 VSS.n6165 VSS.n6164 0.13
R20653 VSS.n6173 VSS.n6172 0.13
R20654 VSS.n6181 VSS.n6180 0.13
R20655 VSS.n6244 VSS.n6188 0.13
R20656 VSS.n10550 VSS.n10549 0.119
R20657 VSS.n17764 VSS.n17763 0.116
R20658 VSS.n18021 VSS 0.108
R20659 VSS.n16588 VSS.n16587 0.101
R20660 VSS.n12637 VSS.n12636 0.101
R20661 VSS.n9205 VSS.n9204 0.101
R20662 VSS.t171 VSS.t176 0.101
R20663 VSS.t162 VSS.t164 0.101
R20664 VSS.t179 VSS.t170 0.101
R20665 VSS.t161 VSS.t173 0.101
R20666 VSS.t168 VSS.t174 0.101
R20667 VSS.t166 VSS.t178 0.101
R20668 VSS.t211 VSS.t216 0.101
R20669 VSS.t202 VSS.t204 0.101
R20670 VSS.t219 VSS.t210 0.101
R20671 VSS.t201 VSS.t213 0.101
R20672 VSS.t208 VSS.t214 0.101
R20673 VSS.t206 VSS.t218 0.101
R20674 VSS.t209 VSS.t203 0.101
R20675 VSS.t217 VSS.t205 0.101
R20676 VSS.t215 VSS.t207 0.101
R20677 VSS.t212 VSS.t200 0.101
R20678 VSS.t160 VSS.t172 0.101
R20679 VSS.t175 VSS.t167 0.101
R20680 VSS.t177 VSS.t165 0.101
R20681 VSS.t169 VSS.t163 0.101
R20682 VSS.t191 VSS.t196 0.101
R20683 VSS.t182 VSS.t184 0.101
R20684 VSS.t199 VSS.t190 0.101
R20685 VSS.t181 VSS.t193 0.101
R20686 VSS.t188 VSS.t194 0.101
R20687 VSS.t186 VSS.t198 0.101
R20688 VSS.t189 VSS.t183 0.101
R20689 VSS.t180 VSS.t192 0.101
R20690 VSS.t195 VSS.t187 0.101
R20691 VSS.t197 VSS.t185 0.101
R20692 VSS.t131 VSS.t136 0.101
R20693 VSS.t122 VSS.t124 0.101
R20694 VSS.t140 VSS.t152 0.101
R20695 VSS.t155 VSS.t147 0.101
R20696 VSS.t157 VSS.t145 0.101
R20697 VSS.t149 VSS.t143 0.101
R20698 VSS.t146 VSS.t158 0.101
R20699 VSS.t148 VSS.t154 0.101
R20700 VSS.t141 VSS.t153 0.101
R20701 VSS.t159 VSS.t150 0.101
R20702 VSS.t142 VSS.t144 0.101
R20703 VSS.t151 VSS.t156 0.101
R20704 VSS.t120 VSS.t132 0.101
R20705 VSS.t135 VSS.t127 0.101
R20706 VSS.t137 VSS.t125 0.101
R20707 VSS.t129 VSS.t123 0.101
R20708 VSS.t126 VSS.t138 0.101
R20709 VSS.t128 VSS.t134 0.101
R20710 VSS.t121 VSS.t133 0.101
R20711 VSS.t139 VSS.t130 0.101
R20712 VSS.n17765 VSS.n17764 0.096
R20713 VSS.n7045 VSS.n7044 0.091
R20714 VSS.n437 VSS.n343 0.089
R20715 VSS.n5784 VSS.n5783 0.087
R20716 VSS.n18022 VSS 0.079
R20717 VSS.n18025 VSS 0.079
R20718 VSS.n0  0.077
R20719  VSS.n18327 0.077
R20720 VSS.n286 VSS.n285 0.077
R20721 VSS.n23 VSS.n18 0.077
R20722 VSS.n17623 VSS.n17618 0.077
R20723 VSS.n14113 VSS.n14108 0.077
R20724 VSS.n10591 VSS.n10586 0.077
R20725 VSS.n7073 VSS.n7068 0.077
R20726 VSS.n510 VSS.n505 0.077
R20727 VSS.n452 VSS.n447 0.077
R20728 VSS.n313 VSS.n308 0.077
R20729 VSS.n302 VSS.n297 0.077
R20730 VSS.n18118 VSS.n18113 0.077
R20731 VSS.n18256 VSS.n18255 0.077
R20732 VSS.n18321 VSS.n18320 0.076
R20733 VSS.n221 VSS.n216 0.076
R20734 VSS.n50 VSS.n49 0.076
R20735 VSS.n69 VSS.n68 0.076
R20736 VSS.n90 VSS.n89 0.076
R20737 VSS.n111 VSS.n110 0.076
R20738 VSS.n132 VSS.n131 0.076
R20739 VSS.n153 VSS.n152 0.076
R20740 VSS.n174 VSS.n173 0.076
R20741 VSS.n195 VSS.n194 0.076
R20742 VSS.n250 VSS.n245 0.076
R20743 VSS.n18273 VSS.n18272 0.076
R20744 VSS.n271 VSS.n270 0.074
R20745 VSS.n237 VSS.n236 0.074
R20746 VSS.n18090 VSS.n31 0.074
R20747 VSS.n18089 VSS.n32 0.074
R20748 VSS.n17643 VSS.n17631 0.074
R20749 VSS.n17642 VSS.n17632 0.074
R20750 VSS.n17611 VSS.n14120 0.074
R20751 VSS.n17609 VSS.n17599 0.074
R20752 VSS.n14101 VSS.n10599 0.074
R20753 VSS.n14095 VSS.n14085 0.074
R20754 VSS.n10579 VSS.n7080 0.074
R20755 VSS.n10577 VSS.n10567 0.074
R20756 VSS.n7061 VSS.n517 0.074
R20757 VSS.n7058 VSS.n7048 0.074
R20758 VSS.n498 VSS.n459 0.074
R20759 VSS.n470 VSS.n460 0.074
R20760 VSS.n440 VSS.n321 0.074
R20761 VSS.n342 VSS.n332 0.074
R20762 VSS.n17741 VSS.n17740 0.074
R20763 VSS.n18027 VSS.n257 0.074
R20764 VSS.n18134 VSS.n18133 0.074
R20765 VSS.n18295 VSS.n18294 0.074
R20766 VSS.n16571 VSS 0.066
R20767 VSS.n12620 VSS 0.066
R20768 VSS.n9188 VSS 0.066
R20769 VSS.n5131 VSS.n5130 0.066
R20770 VSS.n3094 VSS.n3093 0.066
R20771 VSS.n1168 VSS 0.066
R20772 VSS.n6189 VSS 0.066
R20773 VSS.n17764 VSS.n17761 0.062
R20774 VSS.n18026 VSS 0.056
R20775 VSS.n16589 VSS 0.053
R20776 VSS.n9206 VSS 0.053
R20777 VSS.n14082 VSS.n10600 0.051
R20778 VSS.n18327 VSS 0.05
R20779 VSS.n260  0.05
R20780 VSS.n7047 VSS.n518 0.048
R20781 VSS.n495 VSS.n493 0.043
R20782 VSS.n5784 VSS.n519 0.042
R20783 VSS.n18234 VSS.n18233 0.042
R20784 VSS.n18292 VSS.n18291 0.042
R20785 VSS.n18235 VSS.n12 0.041
R20786 VSS.n18290 VSS.n18289 0.041
R20787 VSS.n400 VSS.n399 0.04
R20788 VSS.n416 VSS.n355 0.04
R20789 VSS.n18192 VSS.n18191 0.04
R20790 VSS.n18208 VSS.n18147 0.04
R20791 VSS.n10566 VSS.n7082 0.038
R20792 VSS.n12 VSS.n11 0.036
R20793 VSS.n18289 VSS.n18288 0.036
R20794 VSS.n18233 VSS.n18232 0.036
R20795 VSS.n18293 VSS.n18292 0.036
R20796 VSS.n17753 VSS.n17752 0.036
R20797 VSS.n389 VSS.n364 0.035
R20798 VSS.n423 VSS.n351 0.035
R20799 VSS.n18181 VSS.n18156 0.035
R20800 VSS.n18209 VSS.n18141 0.035
R20801 VSS.n259  0.033
R20802 VSS.n260  0.033
R20803 VSS.n14081 VSS.n14080 0.032
R20804 VSS.n492 VSS.n491 0.029
R20805 VSS.n382 VSS.n369 0.029
R20806 VSS.n431 VSS.n346 0.029
R20807 VSS.n18174 VSS.n18161 0.029
R20808 VSS.n18219 VSS.n18218 0.029
R20809 VSS.n16588 VSS.n16526 0.028
R20810 VSS.n12637 VSS.n12575 0.028
R20811 VSS.n9205 VSS.n9143 0.028
R20812 VSS.n331 VSS.n330 0.028
R20813 VSS.n10564 VSS.n10550 0.027
R20814 VSS.n7046 VSS.n7045 0.025
R20815 VSS.n376 VSS.n373 0.024
R20816 VSS.n433 VSS.n343 0.024
R20817 VSS.n18168 VSS.n18165 0.024
R20818 VSS.n18228 VSS.n18136 0.024
R20819 VSS.n18038 VSS.n18037 0.024
R20820 VSS.n18040 VSS.n18039 0.024
R20821 VSS.n18303 VSS.n18300 0.024
R20822 VSS.n18126 VSS.n18125 0.024
R20823 VSS.n18124 VSS.n18123 0.024
R20824 VSS.n0  0.023
R20825 VSS.n259  0.023
R20826 VSS.n10565 VSS.n7084 0.023
R20827 VSS.n486 VSS.t171 0.023
R20828 VSS.n487 VSS.t162 0.023
R20829 VSS.n488 VSS.t179 0.023
R20830 VSS.n489 VSS.t161 0.023
R20831 VSS.n490 VSS.t168 0.023
R20832 VSS.n491 VSS.t166 0.023
R20833 VSS.n473 VSS.t211 0.023
R20834 VSS.n474 VSS.t202 0.023
R20835 VSS.n475 VSS.t219 0.023
R20836 VSS.n476 VSS.t201 0.023
R20837 VSS.n477 VSS.t208 0.023
R20838 VSS.n478 VSS.t206 0.023
R20839 VSS.n479 VSS.t209 0.023
R20840 VSS.n480 VSS.t217 0.023
R20841 VSS.n481 VSS.t215 0.023
R20842 VSS.n482 VSS.t160 0.023
R20843 VSS.n483 VSS.t175 0.023
R20844 VSS.n484 VSS.t177 0.023
R20845 VSS.n485 VSS.t169 0.023
R20846 VSS.n322 VSS.t191 0.023
R20847 VSS.n323 VSS.t182 0.023
R20848 VSS.n324 VSS.t199 0.023
R20849 VSS.n325 VSS.t181 0.023
R20850 VSS.n326 VSS.t188 0.023
R20851 VSS.n327 VSS.t186 0.023
R20852 VSS.n328 VSS.t189 0.023
R20853 VSS.n329 VSS.t195 0.023
R20854 VSS.n330 VSS.t197 0.023
R20855 VSS.n17762 VSS.t131 0.023
R20856 VSS.n17763 VSS.t122 0.023
R20857 VSS.n17744 VSS.t155 0.023
R20858 VSS.n17745 VSS.t157 0.023
R20859 VSS.n17746 VSS.t149 0.023
R20860 VSS.n17747 VSS.t146 0.023
R20861 VSS.n17748 VSS.t148 0.023
R20862 VSS.n17749 VSS.t141 0.023
R20863 VSS.n17750 VSS.t159 0.023
R20864 VSS.n17751 VSS.t142 0.023
R20865 VSS.n17752 VSS.t151 0.023
R20866 VSS.n17754 VSS.t120 0.023
R20867 VSS.n17755 VSS.t135 0.023
R20868 VSS.n17756 VSS.t137 0.023
R20869 VSS.n17757 VSS.t129 0.023
R20870 VSS.n17758 VSS.t126 0.023
R20871 VSS.n17759 VSS.t128 0.023
R20872 VSS.n17760 VSS.t121 0.023
R20873 VSS.n17761 VSS.t139 0.023
R20874 VSS.n18257 VSS.n18256 0.023
R20875 VSS.n6938 VSS.n5785 0.022
R20876 VSS.n265 VSS.n264 0.021
R20877 VSS.n289 VSS.n288 0.021
R20878 VSS.n225 VSS.n223 0.021
R20879 VSS.n231 VSS.n230 0.021
R20880 VSS.n209 VSS.n208 0.021
R20881 VSS.n18086 VSS.n18085 0.021
R20882 VSS.n17639 VSS.n17638 0.021
R20883 VSS.n17606 VSS.n17605 0.021
R20884 VSS.n14092 VSS.n14091 0.021
R20885 VSS.n10574 VSS.n10573 0.021
R20886 VSS.n7055 VSS.n7054 0.021
R20887 VSS.n467 VSS.n466 0.021
R20888 VSS.n339 VSS.n338 0.021
R20889 VSS.n52 VSS.n44 0.021
R20890 VSS.n43 VSS.n41 0.021
R20891 VSS.n18086 VSS.n37 0.021
R20892 VSS.n71 VSS.n63 0.021
R20893 VSS.n62 VSS.n60 0.021
R20894 VSS.n17639 VSS.n17637 0.021
R20895 VSS.n92 VSS.n84 0.021
R20896 VSS.n83 VSS.n81 0.021
R20897 VSS.n17606 VSS.n17604 0.021
R20898 VSS.n113 VSS.n105 0.021
R20899 VSS.n104 VSS.n102 0.021
R20900 VSS.n14092 VSS.n14090 0.021
R20901 VSS.n134 VSS.n126 0.021
R20902 VSS.n125 VSS.n123 0.021
R20903 VSS.n10574 VSS.n10572 0.021
R20904 VSS.n155 VSS.n147 0.021
R20905 VSS.n146 VSS.n144 0.021
R20906 VSS.n7055 VSS.n7053 0.021
R20907 VSS.n176 VSS.n168 0.021
R20908 VSS.n167 VSS.n165 0.021
R20909 VSS.n467 VSS.n465 0.021
R20910 VSS.n197 VSS.n189 0.021
R20911 VSS.n188 VSS.n186 0.021
R20912 VSS.n339 VSS.n337 0.021
R20913 VSS.n225 VSS.n224 0.021
R20914 VSS.n239 VSS.n235 0.021
R20915 VSS.n14080 VSS.n14079 0.021
R20916 VSS.n381 VSS.n373 0.021
R20917 VSS.n433 VSS.n432 0.021
R20918 VSS.n18173 VSS.n18165 0.021
R20919 VSS.n18138 VSS.n18136 0.021
R20920 VSS.n249 VSS.n248 0.021
R20921 VSS.n17665 VSS.n17664 0.021
R20922 VSS.n17686 VSS.n17685 0.021
R20923 VSS.n17697 VSS.n17696 0.021
R20924 VSS.n17708 VSS.n17707 0.021
R20925 VSS.n28 VSS.n27 0.021
R20926 VSS.n17628 VSS.n17627 0.021
R20927 VSS.n10596 VSS.n10595 0.021
R20928 VSS.n318 VSS.n317 0.021
R20929 VSS.n278 VSS.n276 0.021
R20930 VSS.n284 VSS.n283 0.021
R20931 VSS.n36 VSS.n35 0.021
R20932 VSS.n17636 VSS.n17635 0.021
R20933 VSS.n17603 VSS.n17602 0.021
R20934 VSS.n14089 VSS.n14088 0.021
R20935 VSS.n10571 VSS.n10570 0.021
R20936 VSS.n7052 VSS.n7051 0.021
R20937 VSS.n464 VSS.n463 0.021
R20938 VSS.n336 VSS.n335 0.021
R20939 VSS.n18041 VSS.n254 0.019
R20940 VSS.n18128 VSS.n18127 0.019
R20941 VSS.n17766 VSS.n17742 0.019
R20942 VSS.n18094 VSS.n18093 0.018
R20943 VSS.n17647 VSS.n17646 0.018
R20944 VSS.n17615 VSS.n17614 0.018
R20945 VSS.n14105 VSS.n14104 0.018
R20946 VSS.n10583 VSS.n10582 0.018
R20947 VSS.n7065 VSS.n7064 0.018
R20948 VSS.n502 VSS.n501 0.018
R20949 VSS.n444 VSS.n443 0.018
R20950 VSS.n17738 VSS.n17737 0.018
R20951 VSS.n18031 VSS.n18030 0.018
R20952 VSS.n16 VSS.n15 0.018
R20953 VSS.n18117 VSS.n18116 0.018
R20954 VSS.n18299 VSS.n18298 0.018
R20955 VSS.n18287 VSS.n18286 0.018
R20956 VSS.n18284 VSS.n18283 0.018
R20957 VSS.n18279 VSS.n18278 0.018
R20958 VSS.n18274 VSS.n18273 0.018
R20959 VSS.n14659 VSS.n14644 0.017
R20960 VSS.n14673 VSS.n14661 0.017
R20961 VSS.n14687 VSS.n14675 0.017
R20962 VSS.n14701 VSS.n14689 0.017
R20963 VSS.n14715 VSS.n14703 0.017
R20964 VSS.n14734 VSS.n14717 0.017
R20965 VSS.n14738 VSS.n14737 0.017
R20966 VSS.n14751 VSS.n14594 0.017
R20967 VSS.n14765 VSS.n14753 0.017
R20968 VSS.n14779 VSS.n14767 0.017
R20969 VSS.n14793 VSS.n14781 0.017
R20970 VSS.n14810 VSS.n14795 0.017
R20971 VSS.n14915 VSS.n14903 0.017
R20972 VSS.n14929 VSS.n14917 0.017
R20973 VSS.n14943 VSS.n14931 0.017
R20974 VSS.n14957 VSS.n14945 0.017
R20975 VSS.n14971 VSS.n14959 0.017
R20976 VSS.n14990 VSS.n14973 0.017
R20977 VSS.n14994 VSS.n14993 0.017
R20978 VSS.n15007 VSS.n14588 0.017
R20979 VSS.n15021 VSS.n15009 0.017
R20980 VSS.n15035 VSS.n15023 0.017
R20981 VSS.n15049 VSS.n15037 0.017
R20982 VSS.n15066 VSS.n15051 0.017
R20983 VSS.n15159 VSS.n15147 0.017
R20984 VSS.n15173 VSS.n15161 0.017
R20985 VSS.n15187 VSS.n15175 0.017
R20986 VSS.n15201 VSS.n15189 0.017
R20987 VSS.n15215 VSS.n15203 0.017
R20988 VSS.n15234 VSS.n15217 0.017
R20989 VSS.n15238 VSS.n15237 0.017
R20990 VSS.n15251 VSS.n14582 0.017
R20991 VSS.n15265 VSS.n15253 0.017
R20992 VSS.n15279 VSS.n15267 0.017
R20993 VSS.n15293 VSS.n15281 0.017
R20994 VSS.n15310 VSS.n15295 0.017
R20995 VSS.n15403 VSS.n15391 0.017
R20996 VSS.n15417 VSS.n15405 0.017
R20997 VSS.n15431 VSS.n15419 0.017
R20998 VSS.n15445 VSS.n15433 0.017
R20999 VSS.n15459 VSS.n15447 0.017
R21000 VSS.n15478 VSS.n15461 0.017
R21001 VSS.n15482 VSS.n15481 0.017
R21002 VSS.n15495 VSS.n14576 0.017
R21003 VSS.n15509 VSS.n15497 0.017
R21004 VSS.n15523 VSS.n15511 0.017
R21005 VSS.n15537 VSS.n15525 0.017
R21006 VSS.n15554 VSS.n15539 0.017
R21007 VSS.n15647 VSS.n15635 0.017
R21008 VSS.n15661 VSS.n15649 0.017
R21009 VSS.n15675 VSS.n15663 0.017
R21010 VSS.n15689 VSS.n15677 0.017
R21011 VSS.n15703 VSS.n15691 0.017
R21012 VSS.n15722 VSS.n15705 0.017
R21013 VSS.n15726 VSS.n15725 0.017
R21014 VSS.n15739 VSS.n14570 0.017
R21015 VSS.n15753 VSS.n15741 0.017
R21016 VSS.n15767 VSS.n15755 0.017
R21017 VSS.n15781 VSS.n15769 0.017
R21018 VSS.n15798 VSS.n15783 0.017
R21019 VSS.n15891 VSS.n15879 0.017
R21020 VSS.n15905 VSS.n15893 0.017
R21021 VSS.n15919 VSS.n15907 0.017
R21022 VSS.n15933 VSS.n15921 0.017
R21023 VSS.n15947 VSS.n15935 0.017
R21024 VSS.n15966 VSS.n15949 0.017
R21025 VSS.n15970 VSS.n15969 0.017
R21026 VSS.n15983 VSS.n14564 0.017
R21027 VSS.n15997 VSS.n15985 0.017
R21028 VSS.n16011 VSS.n15999 0.017
R21029 VSS.n16025 VSS.n16013 0.017
R21030 VSS.n16042 VSS.n16027 0.017
R21031 VSS.n16135 VSS.n16123 0.017
R21032 VSS.n16149 VSS.n16137 0.017
R21033 VSS.n16163 VSS.n16151 0.017
R21034 VSS.n16177 VSS.n16165 0.017
R21035 VSS.n16191 VSS.n16179 0.017
R21036 VSS.n16210 VSS.n16193 0.017
R21037 VSS.n16214 VSS.n16213 0.017
R21038 VSS.n16227 VSS.n14558 0.017
R21039 VSS.n16241 VSS.n16229 0.017
R21040 VSS.n16255 VSS.n16243 0.017
R21041 VSS.n16269 VSS.n16257 0.017
R21042 VSS.n16286 VSS.n16271 0.017
R21043 VSS.n16391 VSS.n16379 0.017
R21044 VSS.n16405 VSS.n16393 0.017
R21045 VSS.n16419 VSS.n16407 0.017
R21046 VSS.n16433 VSS.n16421 0.017
R21047 VSS.n16447 VSS.n16435 0.017
R21048 VSS.n16466 VSS.n16449 0.017
R21049 VSS.n16470 VSS.n16469 0.017
R21050 VSS.n16483 VSS.n14552 0.017
R21051 VSS.n16497 VSS.n16485 0.017
R21052 VSS.n16511 VSS.n16499 0.017
R21053 VSS.n16525 VSS.n16513 0.017
R21054 VSS.n16587 VSS.n16586 0.017
R21055 VSS.n14143 VSS.n14133 0.017
R21056 VSS.n14155 VSS.n14145 0.017
R21057 VSS.n14167 VSS.n14157 0.017
R21058 VSS.n14179 VSS.n14169 0.017
R21059 VSS.n14191 VSS.n14181 0.017
R21060 VSS.n14203 VSS.n14193 0.017
R21061 VSS.n14215 VSS.n14205 0.017
R21062 VSS.n14227 VSS.n14217 0.017
R21063 VSS.n14284 VSS.n14229 0.017
R21064 VSS.n14323 VSS.n14313 0.017
R21065 VSS.n14335 VSS.n14325 0.017
R21066 VSS.n14347 VSS.n14337 0.017
R21067 VSS.n14359 VSS.n14349 0.017
R21068 VSS.n14371 VSS.n14361 0.017
R21069 VSS.n14383 VSS.n14373 0.017
R21070 VSS.n14395 VSS.n14385 0.017
R21071 VSS.n14407 VSS.n14397 0.017
R21072 VSS.n14464 VSS.n14409 0.017
R21073 VSS.n17585 VSS.n17584 0.017
R21074 VSS.n17526 VSS.n17525 0.017
R21075 VSS.n17514 VSS.n17513 0.017
R21076 VSS.n17502 VSS.n17501 0.017
R21077 VSS.n17490 VSS.n17489 0.017
R21078 VSS.n17478 VSS.n17468 0.017
R21079 VSS.n17466 VSS.n17465 0.017
R21080 VSS.n17454 VSS.n17453 0.017
R21081 VSS.n17442 VSS.n17441 0.017
R21082 VSS.n17417 VSS.n17416 0.017
R21083 VSS.n17358 VSS.n17357 0.017
R21084 VSS.n17346 VSS.n17345 0.017
R21085 VSS.n17334 VSS.n17333 0.017
R21086 VSS.n17322 VSS.n17321 0.017
R21087 VSS.n17310 VSS.n17300 0.017
R21088 VSS.n17298 VSS.n17297 0.017
R21089 VSS.n17286 VSS.n17285 0.017
R21090 VSS.n17274 VSS.n17273 0.017
R21091 VSS.n17249 VSS.n17248 0.017
R21092 VSS.n17190 VSS.n17189 0.017
R21093 VSS.n17178 VSS.n17177 0.017
R21094 VSS.n17166 VSS.n17165 0.017
R21095 VSS.n17154 VSS.n17153 0.017
R21096 VSS.n17142 VSS.n17132 0.017
R21097 VSS.n17130 VSS.n17129 0.017
R21098 VSS.n17118 VSS.n17117 0.017
R21099 VSS.n17106 VSS.n17105 0.017
R21100 VSS.n17081 VSS.n17080 0.017
R21101 VSS.n17022 VSS.n17021 0.017
R21102 VSS.n17010 VSS.n17009 0.017
R21103 VSS.n16998 VSS.n16997 0.017
R21104 VSS.n16986 VSS.n16985 0.017
R21105 VSS.n16974 VSS.n16964 0.017
R21106 VSS.n16962 VSS.n16961 0.017
R21107 VSS.n16950 VSS.n16949 0.017
R21108 VSS.n16938 VSS.n16937 0.017
R21109 VSS.n16913 VSS.n16912 0.017
R21110 VSS.n16854 VSS.n16853 0.017
R21111 VSS.n16842 VSS.n16841 0.017
R21112 VSS.n16830 VSS.n16829 0.017
R21113 VSS.n16818 VSS.n16817 0.017
R21114 VSS.n16806 VSS.n16796 0.017
R21115 VSS.n16794 VSS.n16793 0.017
R21116 VSS.n16782 VSS.n16781 0.017
R21117 VSS.n16770 VSS.n16769 0.017
R21118 VSS.n16745 VSS.n16744 0.017
R21119 VSS.n16686 VSS.n16685 0.017
R21120 VSS.n16674 VSS.n16673 0.017
R21121 VSS.n16662 VSS.n16661 0.017
R21122 VSS.n16650 VSS.n16649 0.017
R21123 VSS.n16638 VSS.n16628 0.017
R21124 VSS.n16626 VSS.n16625 0.017
R21125 VSS.n16614 VSS.n16613 0.017
R21126 VSS.n16602 VSS.n16601 0.017
R21127 VSS.n10708 VSS.n10693 0.017
R21128 VSS.n10722 VSS.n10710 0.017
R21129 VSS.n10736 VSS.n10724 0.017
R21130 VSS.n10750 VSS.n10738 0.017
R21131 VSS.n10764 VSS.n10752 0.017
R21132 VSS.n10783 VSS.n10766 0.017
R21133 VSS.n10787 VSS.n10786 0.017
R21134 VSS.n10800 VSS.n10643 0.017
R21135 VSS.n10814 VSS.n10802 0.017
R21136 VSS.n10828 VSS.n10816 0.017
R21137 VSS.n10842 VSS.n10830 0.017
R21138 VSS.n10859 VSS.n10844 0.017
R21139 VSS.n10964 VSS.n10952 0.017
R21140 VSS.n10978 VSS.n10966 0.017
R21141 VSS.n10992 VSS.n10980 0.017
R21142 VSS.n11006 VSS.n10994 0.017
R21143 VSS.n11020 VSS.n11008 0.017
R21144 VSS.n11039 VSS.n11022 0.017
R21145 VSS.n11043 VSS.n11042 0.017
R21146 VSS.n11056 VSS.n10637 0.017
R21147 VSS.n11070 VSS.n11058 0.017
R21148 VSS.n11084 VSS.n11072 0.017
R21149 VSS.n11098 VSS.n11086 0.017
R21150 VSS.n11115 VSS.n11100 0.017
R21151 VSS.n11208 VSS.n11196 0.017
R21152 VSS.n11222 VSS.n11210 0.017
R21153 VSS.n11236 VSS.n11224 0.017
R21154 VSS.n11250 VSS.n11238 0.017
R21155 VSS.n11264 VSS.n11252 0.017
R21156 VSS.n11283 VSS.n11266 0.017
R21157 VSS.n11287 VSS.n11286 0.017
R21158 VSS.n11300 VSS.n10631 0.017
R21159 VSS.n11314 VSS.n11302 0.017
R21160 VSS.n11328 VSS.n11316 0.017
R21161 VSS.n11342 VSS.n11330 0.017
R21162 VSS.n11359 VSS.n11344 0.017
R21163 VSS.n11452 VSS.n11440 0.017
R21164 VSS.n11466 VSS.n11454 0.017
R21165 VSS.n11480 VSS.n11468 0.017
R21166 VSS.n11494 VSS.n11482 0.017
R21167 VSS.n11508 VSS.n11496 0.017
R21168 VSS.n11527 VSS.n11510 0.017
R21169 VSS.n11531 VSS.n11530 0.017
R21170 VSS.n11544 VSS.n10625 0.017
R21171 VSS.n11558 VSS.n11546 0.017
R21172 VSS.n11572 VSS.n11560 0.017
R21173 VSS.n11586 VSS.n11574 0.017
R21174 VSS.n11603 VSS.n11588 0.017
R21175 VSS.n11696 VSS.n11684 0.017
R21176 VSS.n11710 VSS.n11698 0.017
R21177 VSS.n11724 VSS.n11712 0.017
R21178 VSS.n11738 VSS.n11726 0.017
R21179 VSS.n11752 VSS.n11740 0.017
R21180 VSS.n11771 VSS.n11754 0.017
R21181 VSS.n11775 VSS.n11774 0.017
R21182 VSS.n11788 VSS.n10619 0.017
R21183 VSS.n11802 VSS.n11790 0.017
R21184 VSS.n11816 VSS.n11804 0.017
R21185 VSS.n11830 VSS.n11818 0.017
R21186 VSS.n11847 VSS.n11832 0.017
R21187 VSS.n11940 VSS.n11928 0.017
R21188 VSS.n11954 VSS.n11942 0.017
R21189 VSS.n11968 VSS.n11956 0.017
R21190 VSS.n11982 VSS.n11970 0.017
R21191 VSS.n11996 VSS.n11984 0.017
R21192 VSS.n12015 VSS.n11998 0.017
R21193 VSS.n12019 VSS.n12018 0.017
R21194 VSS.n12032 VSS.n10613 0.017
R21195 VSS.n12046 VSS.n12034 0.017
R21196 VSS.n12060 VSS.n12048 0.017
R21197 VSS.n12074 VSS.n12062 0.017
R21198 VSS.n12091 VSS.n12076 0.017
R21199 VSS.n12184 VSS.n12172 0.017
R21200 VSS.n12198 VSS.n12186 0.017
R21201 VSS.n12212 VSS.n12200 0.017
R21202 VSS.n12226 VSS.n12214 0.017
R21203 VSS.n12240 VSS.n12228 0.017
R21204 VSS.n12259 VSS.n12242 0.017
R21205 VSS.n12263 VSS.n12262 0.017
R21206 VSS.n12276 VSS.n10607 0.017
R21207 VSS.n12290 VSS.n12278 0.017
R21208 VSS.n12304 VSS.n12292 0.017
R21209 VSS.n12318 VSS.n12306 0.017
R21210 VSS.n12335 VSS.n12320 0.017
R21211 VSS.n12440 VSS.n12428 0.017
R21212 VSS.n12454 VSS.n12442 0.017
R21213 VSS.n12468 VSS.n12456 0.017
R21214 VSS.n12482 VSS.n12470 0.017
R21215 VSS.n12496 VSS.n12484 0.017
R21216 VSS.n12515 VSS.n12498 0.017
R21217 VSS.n12519 VSS.n12518 0.017
R21218 VSS.n12532 VSS.n10601 0.017
R21219 VSS.n12546 VSS.n12534 0.017
R21220 VSS.n12560 VSS.n12548 0.017
R21221 VSS.n12574 VSS.n12562 0.017
R21222 VSS.n12636 VSS.n12635 0.017
R21223 VSS.n12660 VSS.n12650 0.017
R21224 VSS.n12672 VSS.n12662 0.017
R21225 VSS.n12684 VSS.n12674 0.017
R21226 VSS.n12696 VSS.n12686 0.017
R21227 VSS.n12708 VSS.n12698 0.017
R21228 VSS.n12720 VSS.n12710 0.017
R21229 VSS.n12732 VSS.n12722 0.017
R21230 VSS.n12744 VSS.n12734 0.017
R21231 VSS.n12801 VSS.n12746 0.017
R21232 VSS.n12840 VSS.n12830 0.017
R21233 VSS.n12852 VSS.n12842 0.017
R21234 VSS.n12864 VSS.n12854 0.017
R21235 VSS.n12876 VSS.n12866 0.017
R21236 VSS.n12888 VSS.n12878 0.017
R21237 VSS.n12900 VSS.n12890 0.017
R21238 VSS.n12912 VSS.n12902 0.017
R21239 VSS.n12924 VSS.n12914 0.017
R21240 VSS.n12981 VSS.n12926 0.017
R21241 VSS.n13020 VSS.n13010 0.017
R21242 VSS.n13032 VSS.n13022 0.017
R21243 VSS.n13044 VSS.n13034 0.017
R21244 VSS.n13056 VSS.n13046 0.017
R21245 VSS.n13068 VSS.n13058 0.017
R21246 VSS.n13080 VSS.n13070 0.017
R21247 VSS.n13092 VSS.n13082 0.017
R21248 VSS.n13104 VSS.n13094 0.017
R21249 VSS.n13161 VSS.n13106 0.017
R21250 VSS.n13200 VSS.n13190 0.017
R21251 VSS.n13212 VSS.n13202 0.017
R21252 VSS.n13224 VSS.n13214 0.017
R21253 VSS.n13236 VSS.n13226 0.017
R21254 VSS.n13248 VSS.n13238 0.017
R21255 VSS.n13260 VSS.n13250 0.017
R21256 VSS.n13272 VSS.n13262 0.017
R21257 VSS.n13284 VSS.n13274 0.017
R21258 VSS.n13341 VSS.n13286 0.017
R21259 VSS.n13380 VSS.n13370 0.017
R21260 VSS.n13392 VSS.n13382 0.017
R21261 VSS.n13404 VSS.n13394 0.017
R21262 VSS.n13416 VSS.n13406 0.017
R21263 VSS.n13428 VSS.n13418 0.017
R21264 VSS.n13440 VSS.n13430 0.017
R21265 VSS.n13452 VSS.n13442 0.017
R21266 VSS.n13464 VSS.n13454 0.017
R21267 VSS.n13521 VSS.n13466 0.017
R21268 VSS.n13560 VSS.n13550 0.017
R21269 VSS.n13572 VSS.n13562 0.017
R21270 VSS.n13584 VSS.n13574 0.017
R21271 VSS.n13596 VSS.n13586 0.017
R21272 VSS.n13608 VSS.n13598 0.017
R21273 VSS.n13620 VSS.n13610 0.017
R21274 VSS.n13632 VSS.n13622 0.017
R21275 VSS.n13644 VSS.n13634 0.017
R21276 VSS.n13701 VSS.n13646 0.017
R21277 VSS.n13740 VSS.n13730 0.017
R21278 VSS.n13752 VSS.n13742 0.017
R21279 VSS.n13764 VSS.n13754 0.017
R21280 VSS.n13776 VSS.n13766 0.017
R21281 VSS.n13788 VSS.n13778 0.017
R21282 VSS.n13800 VSS.n13790 0.017
R21283 VSS.n13812 VSS.n13802 0.017
R21284 VSS.n13824 VSS.n13814 0.017
R21285 VSS.n13881 VSS.n13826 0.017
R21286 VSS.n13920 VSS.n13910 0.017
R21287 VSS.n13932 VSS.n13922 0.017
R21288 VSS.n13944 VSS.n13934 0.017
R21289 VSS.n13956 VSS.n13946 0.017
R21290 VSS.n13968 VSS.n13958 0.017
R21291 VSS.n13980 VSS.n13970 0.017
R21292 VSS.n13992 VSS.n13982 0.017
R21293 VSS.n14004 VSS.n13994 0.017
R21294 VSS.n14061 VSS.n14006 0.017
R21295 VSS.n7276 VSS.n7261 0.017
R21296 VSS.n7290 VSS.n7278 0.017
R21297 VSS.n7304 VSS.n7292 0.017
R21298 VSS.n7318 VSS.n7306 0.017
R21299 VSS.n7332 VSS.n7320 0.017
R21300 VSS.n7351 VSS.n7334 0.017
R21301 VSS.n7355 VSS.n7354 0.017
R21302 VSS.n7368 VSS.n7211 0.017
R21303 VSS.n7382 VSS.n7370 0.017
R21304 VSS.n7396 VSS.n7384 0.017
R21305 VSS.n7410 VSS.n7398 0.017
R21306 VSS.n7427 VSS.n7412 0.017
R21307 VSS.n7532 VSS.n7520 0.017
R21308 VSS.n7546 VSS.n7534 0.017
R21309 VSS.n7560 VSS.n7548 0.017
R21310 VSS.n7574 VSS.n7562 0.017
R21311 VSS.n7588 VSS.n7576 0.017
R21312 VSS.n7607 VSS.n7590 0.017
R21313 VSS.n7611 VSS.n7610 0.017
R21314 VSS.n7624 VSS.n7205 0.017
R21315 VSS.n7638 VSS.n7626 0.017
R21316 VSS.n7652 VSS.n7640 0.017
R21317 VSS.n7666 VSS.n7654 0.017
R21318 VSS.n7683 VSS.n7668 0.017
R21319 VSS.n7776 VSS.n7764 0.017
R21320 VSS.n7790 VSS.n7778 0.017
R21321 VSS.n7804 VSS.n7792 0.017
R21322 VSS.n7818 VSS.n7806 0.017
R21323 VSS.n7832 VSS.n7820 0.017
R21324 VSS.n7851 VSS.n7834 0.017
R21325 VSS.n7855 VSS.n7854 0.017
R21326 VSS.n7868 VSS.n7199 0.017
R21327 VSS.n7882 VSS.n7870 0.017
R21328 VSS.n7896 VSS.n7884 0.017
R21329 VSS.n7910 VSS.n7898 0.017
R21330 VSS.n7927 VSS.n7912 0.017
R21331 VSS.n8020 VSS.n8008 0.017
R21332 VSS.n8034 VSS.n8022 0.017
R21333 VSS.n8048 VSS.n8036 0.017
R21334 VSS.n8062 VSS.n8050 0.017
R21335 VSS.n8076 VSS.n8064 0.017
R21336 VSS.n8095 VSS.n8078 0.017
R21337 VSS.n8099 VSS.n8098 0.017
R21338 VSS.n8112 VSS.n7193 0.017
R21339 VSS.n8126 VSS.n8114 0.017
R21340 VSS.n8140 VSS.n8128 0.017
R21341 VSS.n8154 VSS.n8142 0.017
R21342 VSS.n8171 VSS.n8156 0.017
R21343 VSS.n8264 VSS.n8252 0.017
R21344 VSS.n8278 VSS.n8266 0.017
R21345 VSS.n8292 VSS.n8280 0.017
R21346 VSS.n8306 VSS.n8294 0.017
R21347 VSS.n8320 VSS.n8308 0.017
R21348 VSS.n8339 VSS.n8322 0.017
R21349 VSS.n8343 VSS.n8342 0.017
R21350 VSS.n8356 VSS.n7187 0.017
R21351 VSS.n8370 VSS.n8358 0.017
R21352 VSS.n8384 VSS.n8372 0.017
R21353 VSS.n8398 VSS.n8386 0.017
R21354 VSS.n8415 VSS.n8400 0.017
R21355 VSS.n8508 VSS.n8496 0.017
R21356 VSS.n8522 VSS.n8510 0.017
R21357 VSS.n8536 VSS.n8524 0.017
R21358 VSS.n8550 VSS.n8538 0.017
R21359 VSS.n8564 VSS.n8552 0.017
R21360 VSS.n8583 VSS.n8566 0.017
R21361 VSS.n8587 VSS.n8586 0.017
R21362 VSS.n8600 VSS.n7181 0.017
R21363 VSS.n8614 VSS.n8602 0.017
R21364 VSS.n8628 VSS.n8616 0.017
R21365 VSS.n8642 VSS.n8630 0.017
R21366 VSS.n8659 VSS.n8644 0.017
R21367 VSS.n8752 VSS.n8740 0.017
R21368 VSS.n8766 VSS.n8754 0.017
R21369 VSS.n8780 VSS.n8768 0.017
R21370 VSS.n8794 VSS.n8782 0.017
R21371 VSS.n8808 VSS.n8796 0.017
R21372 VSS.n8827 VSS.n8810 0.017
R21373 VSS.n8831 VSS.n8830 0.017
R21374 VSS.n8844 VSS.n7175 0.017
R21375 VSS.n8858 VSS.n8846 0.017
R21376 VSS.n8872 VSS.n8860 0.017
R21377 VSS.n8886 VSS.n8874 0.017
R21378 VSS.n8903 VSS.n8888 0.017
R21379 VSS.n9008 VSS.n8996 0.017
R21380 VSS.n9022 VSS.n9010 0.017
R21381 VSS.n9036 VSS.n9024 0.017
R21382 VSS.n9050 VSS.n9038 0.017
R21383 VSS.n9064 VSS.n9052 0.017
R21384 VSS.n9083 VSS.n9066 0.017
R21385 VSS.n9087 VSS.n9086 0.017
R21386 VSS.n9100 VSS.n7169 0.017
R21387 VSS.n9114 VSS.n9102 0.017
R21388 VSS.n9128 VSS.n9116 0.017
R21389 VSS.n9142 VSS.n9130 0.017
R21390 VSS.n9204 VSS.n9203 0.017
R21391 VSS.n10549 VSS.n10548 0.017
R21392 VSS.n10491 VSS.n10490 0.017
R21393 VSS.n10479 VSS.n10478 0.017
R21394 VSS.n10467 VSS.n10466 0.017
R21395 VSS.n10455 VSS.n10454 0.017
R21396 VSS.n10443 VSS.n10433 0.017
R21397 VSS.n10431 VSS.n10430 0.017
R21398 VSS.n10419 VSS.n10418 0.017
R21399 VSS.n10407 VSS.n10406 0.017
R21400 VSS.n10381 VSS.n10380 0.017
R21401 VSS.n10324 VSS.n10323 0.017
R21402 VSS.n10312 VSS.n10311 0.017
R21403 VSS.n10300 VSS.n10299 0.017
R21404 VSS.n10288 VSS.n10287 0.017
R21405 VSS.n10276 VSS.n10266 0.017
R21406 VSS.n10264 VSS.n10263 0.017
R21407 VSS.n10252 VSS.n10251 0.017
R21408 VSS.n10240 VSS.n10239 0.017
R21409 VSS.n10213 VSS.n10212 0.017
R21410 VSS.n10156 VSS.n10155 0.017
R21411 VSS.n10144 VSS.n10143 0.017
R21412 VSS.n10132 VSS.n10131 0.017
R21413 VSS.n10120 VSS.n10119 0.017
R21414 VSS.n10108 VSS.n10098 0.017
R21415 VSS.n10096 VSS.n10095 0.017
R21416 VSS.n10084 VSS.n10083 0.017
R21417 VSS.n10072 VSS.n10071 0.017
R21418 VSS.n10045 VSS.n10044 0.017
R21419 VSS.n9988 VSS.n9987 0.017
R21420 VSS.n9976 VSS.n9975 0.017
R21421 VSS.n9964 VSS.n9963 0.017
R21422 VSS.n9952 VSS.n9951 0.017
R21423 VSS.n9940 VSS.n9930 0.017
R21424 VSS.n9928 VSS.n9927 0.017
R21425 VSS.n9916 VSS.n9915 0.017
R21426 VSS.n9904 VSS.n9903 0.017
R21427 VSS.n9877 VSS.n9876 0.017
R21428 VSS.n9820 VSS.n9819 0.017
R21429 VSS.n9808 VSS.n9807 0.017
R21430 VSS.n9796 VSS.n9795 0.017
R21431 VSS.n9784 VSS.n9783 0.017
R21432 VSS.n9772 VSS.n9762 0.017
R21433 VSS.n9760 VSS.n9759 0.017
R21434 VSS.n9748 VSS.n9747 0.017
R21435 VSS.n9736 VSS.n9735 0.017
R21436 VSS.n9709 VSS.n9708 0.017
R21437 VSS.n9652 VSS.n9651 0.017
R21438 VSS.n9640 VSS.n9639 0.017
R21439 VSS.n9628 VSS.n9627 0.017
R21440 VSS.n9616 VSS.n9615 0.017
R21441 VSS.n9604 VSS.n9594 0.017
R21442 VSS.n9592 VSS.n9591 0.017
R21443 VSS.n9580 VSS.n9579 0.017
R21444 VSS.n9568 VSS.n9567 0.017
R21445 VSS.n9541 VSS.n9540 0.017
R21446 VSS.n9484 VSS.n9483 0.017
R21447 VSS.n9472 VSS.n9471 0.017
R21448 VSS.n9460 VSS.n9459 0.017
R21449 VSS.n9448 VSS.n9447 0.017
R21450 VSS.n9436 VSS.n9426 0.017
R21451 VSS.n9424 VSS.n9423 0.017
R21452 VSS.n9412 VSS.n9411 0.017
R21453 VSS.n9400 VSS.n9399 0.017
R21454 VSS.n9373 VSS.n9372 0.017
R21455 VSS.n9316 VSS.n9315 0.017
R21456 VSS.n9304 VSS.n9303 0.017
R21457 VSS.n9292 VSS.n9291 0.017
R21458 VSS.n9280 VSS.n9279 0.017
R21459 VSS.n9268 VSS.n9258 0.017
R21460 VSS.n9256 VSS.n9255 0.017
R21461 VSS.n9244 VSS.n9243 0.017
R21462 VSS.n9232 VSS.n9231 0.017
R21463 VSS.n3459 VSS.n3453 0.017
R21464 VSS.n3798 VSS.n3797 0.017
R21465 VSS.n3786 VSS.n3462 0.017
R21466 VSS.n3784 VSS.n3468 0.017
R21467 VSS.n3775 VSS.n3774 0.017
R21468 VSS.n3763 VSS.n3481 0.017
R21469 VSS.n3761 VSS.n3487 0.017
R21470 VSS.n3752 VSS.n3751 0.017
R21471 VSS.n3740 VSS.n3500 0.017
R21472 VSS.n3738 VSS.n3506 0.017
R21473 VSS.n3729 VSS.n3728 0.017
R21474 VSS.n3717 VSS.n3519 0.017
R21475 VSS.n3714 VSS.n3559 0.017
R21476 VSS.n3705 VSS.n3704 0.017
R21477 VSS.n3693 VSS.n3574 0.017
R21478 VSS.n3691 VSS.n3580 0.017
R21479 VSS.n3682 VSS.n3681 0.017
R21480 VSS.n3670 VSS.n3593 0.017
R21481 VSS.n3668 VSS.n3599 0.017
R21482 VSS.n3659 VSS.n3658 0.017
R21483 VSS.n3647 VSS.n3612 0.017
R21484 VSS.n3645 VSS.n3618 0.017
R21485 VSS.n3636 VSS.n3635 0.017
R21486 VSS.n3955 VSS.n3954 0.017
R21487 VSS.n3966 VSS.n3965 0.017
R21488 VSS.n3377 VSS.n3375 0.017
R21489 VSS.n3979 VSS.n3369 0.017
R21490 VSS.n3991 VSS.n3990 0.017
R21491 VSS.n4001 VSS.n4000 0.017
R21492 VSS.n3356 VSS.n3354 0.017
R21493 VSS.n4014 VSS.n3348 0.017
R21494 VSS.n4026 VSS.n4025 0.017
R21495 VSS.n4036 VSS.n4035 0.017
R21496 VSS.n3335 VSS.n3333 0.017
R21497 VSS.n4049 VSS.n3327 0.017
R21498 VSS.n4416 VSS.n4415 0.017
R21499 VSS.n4411 VSS.n4060 0.017
R21500 VSS.n4402 VSS.n4401 0.017
R21501 VSS.n4390 VSS.n4074 0.017
R21502 VSS.n4388 VSS.n4080 0.017
R21503 VSS.n4379 VSS.n4378 0.017
R21504 VSS.n4367 VSS.n4093 0.017
R21505 VSS.n4365 VSS.n4099 0.017
R21506 VSS.n4356 VSS.n4355 0.017
R21507 VSS.n4344 VSS.n4112 0.017
R21508 VSS.n4342 VSS.n4118 0.017
R21509 VSS.n4333 VSS.n4332 0.017
R21510 VSS.n4321 VSS.n4131 0.017
R21511 VSS.n4318 VSS.n4171 0.017
R21512 VSS.n4309 VSS.n4308 0.017
R21513 VSS.n4297 VSS.n4186 0.017
R21514 VSS.n4295 VSS.n4192 0.017
R21515 VSS.n4286 VSS.n4285 0.017
R21516 VSS.n4274 VSS.n4205 0.017
R21517 VSS.n4272 VSS.n4211 0.017
R21518 VSS.n4263 VSS.n4262 0.017
R21519 VSS.n4251 VSS.n4224 0.017
R21520 VSS.n4249 VSS.n4230 0.017
R21521 VSS.n4240 VSS.n3222 0.017
R21522 VSS.n4540 VSS.n4539 0.017
R21523 VSS.n4545 VSS.n3213 0.017
R21524 VSS.n4557 VSS.n4556 0.017
R21525 VSS.n4567 VSS.n4566 0.017
R21526 VSS.n3200 VSS.n3198 0.017
R21527 VSS.n4580 VSS.n3192 0.017
R21528 VSS.n4592 VSS.n4591 0.017
R21529 VSS.n4602 VSS.n4601 0.017
R21530 VSS.n3179 VSS.n3177 0.017
R21531 VSS.n4615 VSS.n3171 0.017
R21532 VSS.n4627 VSS.n4626 0.017
R21533 VSS.n4637 VSS.n4636 0.017
R21534 VSS.n4648 VSS.n3157 0.017
R21535 VSS.n5020 VSS.n4650 0.017
R21536 VSS.n5011 VSS.n5010 0.017
R21537 VSS.n4999 VSS.n4664 0.017
R21538 VSS.n4997 VSS.n4670 0.017
R21539 VSS.n4988 VSS.n4987 0.017
R21540 VSS.n4976 VSS.n4683 0.017
R21541 VSS.n4974 VSS.n4689 0.017
R21542 VSS.n4965 VSS.n4964 0.017
R21543 VSS.n4953 VSS.n4702 0.017
R21544 VSS.n4951 VSS.n4708 0.017
R21545 VSS.n4942 VSS.n4941 0.017
R21546 VSS.n4930 VSS.n4721 0.017
R21547 VSS.n4927 VSS.n4761 0.017
R21548 VSS.n4918 VSS.n4917 0.017
R21549 VSS.n4906 VSS.n4776 0.017
R21550 VSS.n4904 VSS.n4782 0.017
R21551 VSS.n4895 VSS.n4894 0.017
R21552 VSS.n4883 VSS.n4795 0.017
R21553 VSS.n4881 VSS.n4801 0.017
R21554 VSS.n4872 VSS.n4871 0.017
R21555 VSS.n4860 VSS.n4814 0.017
R21556 VSS.n4858 VSS.n4820 0.017
R21557 VSS.n4849 VSS.n4848 0.017
R21558 VSS.n4837 VSS.n4833 0.017
R21559 VSS.n2381 VSS.n2326 0.017
R21560 VSS.n2451 VSS.n2450 0.017
R21561 VSS.n2441 VSS.n2383 0.017
R21562 VSS.n2439 VSS.n2385 0.017
R21563 VSS.n2433 VSS.n2391 0.017
R21564 VSS.n2427 VSS.n2395 0.017
R21565 VSS.n2421 VSS.n2398 0.017
R21566 VSS.n2416 VSS.n2401 0.017
R21567 VSS.n2410 VSS.n2404 0.017
R21568 VSS.n2471 VSS.n2236 0.017
R21569 VSS.n2541 VSS.n2540 0.017
R21570 VSS.n2531 VSS.n2473 0.017
R21571 VSS.n2529 VSS.n2475 0.017
R21572 VSS.n2523 VSS.n2481 0.017
R21573 VSS.n2517 VSS.n2485 0.017
R21574 VSS.n2511 VSS.n2488 0.017
R21575 VSS.n2506 VSS.n2491 0.017
R21576 VSS.n2500 VSS.n2494 0.017
R21577 VSS.n2561 VSS.n2146 0.017
R21578 VSS.n2631 VSS.n2630 0.017
R21579 VSS.n2621 VSS.n2563 0.017
R21580 VSS.n2619 VSS.n2565 0.017
R21581 VSS.n2613 VSS.n2571 0.017
R21582 VSS.n2607 VSS.n2575 0.017
R21583 VSS.n2601 VSS.n2578 0.017
R21584 VSS.n2596 VSS.n2581 0.017
R21585 VSS.n2590 VSS.n2584 0.017
R21586 VSS.n2651 VSS.n2056 0.017
R21587 VSS.n2721 VSS.n2720 0.017
R21588 VSS.n2711 VSS.n2653 0.017
R21589 VSS.n2709 VSS.n2655 0.017
R21590 VSS.n2703 VSS.n2661 0.017
R21591 VSS.n2697 VSS.n2665 0.017
R21592 VSS.n2691 VSS.n2668 0.017
R21593 VSS.n2686 VSS.n2671 0.017
R21594 VSS.n2680 VSS.n2674 0.017
R21595 VSS.n2741 VSS.n1966 0.017
R21596 VSS.n2811 VSS.n2810 0.017
R21597 VSS.n2801 VSS.n2743 0.017
R21598 VSS.n2799 VSS.n2745 0.017
R21599 VSS.n2793 VSS.n2751 0.017
R21600 VSS.n2787 VSS.n2755 0.017
R21601 VSS.n2781 VSS.n2758 0.017
R21602 VSS.n2776 VSS.n2761 0.017
R21603 VSS.n2770 VSS.n2764 0.017
R21604 VSS.n2831 VSS.n1876 0.017
R21605 VSS.n2901 VSS.n2900 0.017
R21606 VSS.n2891 VSS.n2833 0.017
R21607 VSS.n2889 VSS.n2835 0.017
R21608 VSS.n2883 VSS.n2841 0.017
R21609 VSS.n2877 VSS.n2845 0.017
R21610 VSS.n2871 VSS.n2848 0.017
R21611 VSS.n2866 VSS.n2851 0.017
R21612 VSS.n2860 VSS.n2854 0.017
R21613 VSS.n2921 VSS.n1786 0.017
R21614 VSS.n2991 VSS.n2990 0.017
R21615 VSS.n2981 VSS.n2923 0.017
R21616 VSS.n2979 VSS.n2925 0.017
R21617 VSS.n2973 VSS.n2931 0.017
R21618 VSS.n2967 VSS.n2935 0.017
R21619 VSS.n2961 VSS.n2938 0.017
R21620 VSS.n2956 VSS.n2941 0.017
R21621 VSS.n2950 VSS.n2944 0.017
R21622 VSS.n3011 VSS.n1696 0.017
R21623 VSS.n3081 VSS.n3080 0.017
R21624 VSS.n3071 VSS.n3013 0.017
R21625 VSS.n3069 VSS.n3015 0.017
R21626 VSS.n3063 VSS.n3021 0.017
R21627 VSS.n3057 VSS.n3025 0.017
R21628 VSS.n3051 VSS.n3028 0.017
R21629 VSS.n3046 VSS.n3031 0.017
R21630 VSS.n3040 VSS.n3034 0.017
R21631 VSS.n1583 VSS.n1581 0.017
R21632 VSS.n5145 VSS.n1575 0.017
R21633 VSS.n5157 VSS.n5156 0.017
R21634 VSS.n5167 VSS.n5166 0.017
R21635 VSS.n1562 VSS.n1560 0.017
R21636 VSS.n5180 VSS.n1554 0.017
R21637 VSS.n5192 VSS.n5191 0.017
R21638 VSS.n5202 VSS.n5201 0.017
R21639 VSS.n1541 VSS.n1539 0.017
R21640 VSS.n5215 VSS.n1531 0.017
R21641 VSS.n5228 VSS.n5227 0.017
R21642 VSS.n5406 VSS.n5405 0.017
R21643 VSS.n5395 VSS.n5394 0.017
R21644 VSS.n5383 VSS.n5238 0.017
R21645 VSS.n5381 VSS.n5245 0.017
R21646 VSS.n5372 VSS.n5371 0.017
R21647 VSS.n5360 VSS.n5258 0.017
R21648 VSS.n5358 VSS.n5264 0.017
R21649 VSS.n5349 VSS.n5348 0.017
R21650 VSS.n5337 VSS.n5277 0.017
R21651 VSS.n5335 VSS.n5283 0.017
R21652 VSS.n5326 VSS.n5325 0.017
R21653 VSS.n5314 VSS.n5296 0.017
R21654 VSS.n5312 VSS.n5303 0.017
R21655 VSS.n1442 VSS.n1440 0.017
R21656 VSS.n5504 VSS.n1434 0.017
R21657 VSS.n5516 VSS.n5515 0.017
R21658 VSS.n5526 VSS.n5525 0.017
R21659 VSS.n1421 VSS.n1419 0.017
R21660 VSS.n5539 VSS.n1413 0.017
R21661 VSS.n5551 VSS.n5550 0.017
R21662 VSS.n5561 VSS.n5560 0.017
R21663 VSS.n1400 VSS.n1398 0.017
R21664 VSS.n5574 VSS.n1390 0.017
R21665 VSS.n5587 VSS.n5586 0.017
R21666 VSS.n5614 VSS.n5613 0.017
R21667 VSS.n5603 VSS.n5602 0.017
R21668 VSS.n5783 VSS.n520 0.017
R21669 VSS.n5774 VSS.n5773 0.017
R21670 VSS.n5762 VSS.n532 0.017
R21671 VSS.n5760 VSS.n538 0.017
R21672 VSS.n5751 VSS.n5750 0.017
R21673 VSS.n5739 VSS.n551 0.017
R21674 VSS.n5737 VSS.n557 0.017
R21675 VSS.n5728 VSS.n5727 0.017
R21676 VSS.n5716 VSS.n570 0.017
R21677 VSS.n5714 VSS.n576 0.017
R21678 VSS.n5705 VSS.n5704 0.017
R21679 VSS.n779 VSS.n777 0.017
R21680 VSS.n790 VSS.n771 0.017
R21681 VSS.n802 VSS.n801 0.017
R21682 VSS.n812 VSS.n811 0.017
R21683 VSS.n758 VSS.n756 0.017
R21684 VSS.n825 VSS.n750 0.017
R21685 VSS.n837 VSS.n836 0.017
R21686 VSS.n847 VSS.n846 0.017
R21687 VSS.n737 VSS.n735 0.017
R21688 VSS.n860 VSS.n729 0.017
R21689 VSS.n872 VSS.n871 0.017
R21690 VSS.n882 VSS.n881 0.017
R21691 VSS.n924 VSS.n923 0.017
R21692 VSS.n707 VSS.n705 0.017
R21693 VSS.n937 VSS.n699 0.017
R21694 VSS.n949 VSS.n948 0.017
R21695 VSS.n959 VSS.n958 0.017
R21696 VSS.n686 VSS.n684 0.017
R21697 VSS.n972 VSS.n678 0.017
R21698 VSS.n984 VSS.n983 0.017
R21699 VSS.n994 VSS.n993 0.017
R21700 VSS.n665 VSS.n663 0.017
R21701 VSS.n1007 VSS.n657 0.017
R21702 VSS.n1265 VSS.n1264 0.017
R21703 VSS.n1260 VSS.n1018 0.017
R21704 VSS.n1251 VSS.n1250 0.017
R21705 VSS.n1239 VSS.n1032 0.017
R21706 VSS.n1237 VSS.n1038 0.017
R21707 VSS.n1228 VSS.n1227 0.017
R21708 VSS.n1216 VSS.n1051 0.017
R21709 VSS.n1214 VSS.n1057 0.017
R21710 VSS.n1205 VSS.n1204 0.017
R21711 VSS.n1193 VSS.n1070 0.017
R21712 VSS.n1191 VSS.n1076 0.017
R21713 VSS.n1182 VSS.n1181 0.017
R21714 VSS.n1170 VSS.n1089 0.017
R21715 VSS.n6675 VSS.n6620 0.017
R21716 VSS.n6744 VSS.n6743 0.017
R21717 VSS.n6734 VSS.n6677 0.017
R21718 VSS.n6732 VSS.n6679 0.017
R21719 VSS.n6726 VSS.n6685 0.017
R21720 VSS.n6720 VSS.n6689 0.017
R21721 VSS.n6714 VSS.n6693 0.017
R21722 VSS.n6708 VSS.n6696 0.017
R21723 VSS.n6703 VSS.n6699 0.017
R21724 VSS.n6765 VSS.n6530 0.017
R21725 VSS.n6834 VSS.n6833 0.017
R21726 VSS.n6824 VSS.n6767 0.017
R21727 VSS.n6822 VSS.n6769 0.017
R21728 VSS.n6816 VSS.n6775 0.017
R21729 VSS.n6810 VSS.n6779 0.017
R21730 VSS.n6804 VSS.n6783 0.017
R21731 VSS.n6798 VSS.n6786 0.017
R21732 VSS.n6793 VSS.n6789 0.017
R21733 VSS.n6855 VSS.n6440 0.017
R21734 VSS.n6924 VSS.n6923 0.017
R21735 VSS.n6914 VSS.n6857 0.017
R21736 VSS.n6912 VSS.n6859 0.017
R21737 VSS.n6906 VSS.n6865 0.017
R21738 VSS.n6900 VSS.n6869 0.017
R21739 VSS.n6894 VSS.n6873 0.017
R21740 VSS.n6888 VSS.n6876 0.017
R21741 VSS.n6883 VSS.n6879 0.017
R21742 VSS.n7044 VSS.n5786 0.017
R21743 VSS.n5798 VSS.n5794 0.017
R21744 VSS.n5804 VSS.n5800 0.017
R21745 VSS.n5810 VSS.n5806 0.017
R21746 VSS.n5815 VSS.n5812 0.017
R21747 VSS.n5822 VSS.n5817 0.017
R21748 VSS.n5828 VSS.n5824 0.017
R21749 VSS.n5834 VSS.n5830 0.017
R21750 VSS.n5839 VSS.n5836 0.017
R21751 VSS.n5893 VSS.n5841 0.017
R21752 VSS.n5901 VSS.n5891 0.017
R21753 VSS.n5909 VSS.n5889 0.017
R21754 VSS.n5917 VSS.n5887 0.017
R21755 VSS.n5925 VSS.n5885 0.017
R21756 VSS.n5933 VSS.n5883 0.017
R21757 VSS.n5941 VSS.n5881 0.017
R21758 VSS.n5949 VSS.n5879 0.017
R21759 VSS.n6372 VSS.n6371 0.017
R21760 VSS.n6009 VSS.n5957 0.017
R21761 VSS.n6017 VSS.n6007 0.017
R21762 VSS.n6025 VSS.n6005 0.017
R21763 VSS.n6033 VSS.n6003 0.017
R21764 VSS.n6041 VSS.n6001 0.017
R21765 VSS.n6049 VSS.n5999 0.017
R21766 VSS.n6057 VSS.n5997 0.017
R21767 VSS.n6065 VSS.n5995 0.017
R21768 VSS.n6308 VSS.n6307 0.017
R21769 VSS.n6125 VSS.n6073 0.017
R21770 VSS.n6133 VSS.n6123 0.017
R21771 VSS.n6141 VSS.n6121 0.017
R21772 VSS.n6149 VSS.n6119 0.017
R21773 VSS.n6157 VSS.n6117 0.017
R21774 VSS.n6165 VSS.n6115 0.017
R21775 VSS.n6173 VSS.n6113 0.017
R21776 VSS.n6181 VSS.n6111 0.017
R21777 VSS.n6244 VSS.n6243 0.017
R21778 VSS.n53 VSS.n52 0.017
R21779 VSS.n59 VSS.n58 0.017
R21780 VSS.n18084 VSS.n18083 0.017
R21781 VSS.n72 VSS.n71 0.017
R21782 VSS.n78 VSS.n77 0.017
R21783 VSS.n80 VSS.n79 0.017
R21784 VSS.n93 VSS.n92 0.017
R21785 VSS.n99 VSS.n98 0.017
R21786 VSS.n101 VSS.n100 0.017
R21787 VSS.n114 VSS.n113 0.017
R21788 VSS.n120 VSS.n119 0.017
R21789 VSS.n122 VSS.n121 0.017
R21790 VSS.n135 VSS.n134 0.017
R21791 VSS.n141 VSS.n140 0.017
R21792 VSS.n143 VSS.n142 0.017
R21793 VSS.n156 VSS.n155 0.017
R21794 VSS.n162 VSS.n161 0.017
R21795 VSS.n164 VSS.n163 0.017
R21796 VSS.n177 VSS.n176 0.017
R21797 VSS.n183 VSS.n182 0.017
R21798 VSS.n185 VSS.n184 0.017
R21799 VSS.n198 VSS.n197 0.017
R21800 VSS.n204 VSS.n203 0.017
R21801 VSS.n206 VSS.n205 0.017
R21802 VSS.n275 VSS.n274 0.017
R21803 VSS.n280 VSS.n279 0.017
R21804 VSS.n291 VSS.n290 0.017
R21805 VSS.n14077 VSS.n14063 0.016
R21806 VSS.n18274 VSS.n18267 0.016
R21807 VSS.n18279 VSS.n18277 0.016
R21808 VSS.n18284 VSS.n18282 0.016
R21809 VSS.n18290 VSS.n18287 0.016
R21810 VSS.n388 VSS.n369 0.016
R21811 VSS.n424 VSS.n346 0.016
R21812 VSS.n18180 VSS.n18161 0.016
R21813 VSS.n18218 VSS.n18217 0.016
R21814 VSS.n275 VSS.n265 0.016
R21815 VSS.n280 VSS.n278 0.016
R21816 VSS.n291 VSS.n289 0.016
R21817 VSS.n53 VSS.n43 0.016
R21818 VSS.n59 VSS.n56 0.016
R21819 VSS.n18086 VSS.n18084 0.016
R21820 VSS.n72 VSS.n62 0.016
R21821 VSS.n78 VSS.n75 0.016
R21822 VSS.n17639 VSS.n80 0.016
R21823 VSS.n93 VSS.n83 0.016
R21824 VSS.n99 VSS.n96 0.016
R21825 VSS.n17606 VSS.n101 0.016
R21826 VSS.n114 VSS.n104 0.016
R21827 VSS.n120 VSS.n117 0.016
R21828 VSS.n14092 VSS.n122 0.016
R21829 VSS.n135 VSS.n125 0.016
R21830 VSS.n141 VSS.n138 0.016
R21831 VSS.n10574 VSS.n143 0.016
R21832 VSS.n156 VSS.n146 0.016
R21833 VSS.n162 VSS.n159 0.016
R21834 VSS.n7055 VSS.n164 0.016
R21835 VSS.n177 VSS.n167 0.016
R21836 VSS.n183 VSS.n180 0.016
R21837 VSS.n467 VSS.n185 0.016
R21838 VSS.n198 VSS.n188 0.016
R21839 VSS.n204 VSS.n201 0.016
R21840 VSS.n339 VSS.n206 0.016
R21841 VSS.n14099 VSS.n14098 0.015
R21842 VSS.n18023 VSS.n18022 0.015
R21843 VSS.n272 VSS.n269 0.015
R21844 VSS.n221 VSS.n220 0.015
R21845 VSS.n18273 VSS.n18271 0.015
R21846 VSS.n18267 VSS.n18265 0.015
R21847 VSS.n18277 VSS.n18275 0.015
R21848 VSS.n18282 VSS.n18280 0.015
R21849 VSS.n18290 VSS.n5 0.015
R21850 VSS.n23 VSS.n22 0.015
R21851 VSS.n50 VSS.n48 0.015
R21852 VSS.n51 VSS.n50 0.015
R21853 VSS.n52 VSS.n51 0.015
R21854 VSS.n43 VSS.n42 0.015
R21855 VSS.n56 VSS.n54 0.015
R21856 VSS.n18087 VSS.n18086 0.015
R21857 VSS.n18088 VSS.n18087 0.015
R21858 VSS.n17623 VSS.n17622 0.015
R21859 VSS.n69 VSS.n67 0.015
R21860 VSS.n70 VSS.n69 0.015
R21861 VSS.n71 VSS.n70 0.015
R21862 VSS.n62 VSS.n61 0.015
R21863 VSS.n75 VSS.n73 0.015
R21864 VSS.n17640 VSS.n17639 0.015
R21865 VSS.n17641 VSS.n17640 0.015
R21866 VSS.n14113 VSS.n14112 0.015
R21867 VSS.n90 VSS.n88 0.015
R21868 VSS.n91 VSS.n90 0.015
R21869 VSS.n92 VSS.n91 0.015
R21870 VSS.n83 VSS.n82 0.015
R21871 VSS.n96 VSS.n94 0.015
R21872 VSS.n17607 VSS.n17606 0.015
R21873 VSS.n17608 VSS.n17607 0.015
R21874 VSS.n10591 VSS.n10590 0.015
R21875 VSS.n111 VSS.n109 0.015
R21876 VSS.n112 VSS.n111 0.015
R21877 VSS.n113 VSS.n112 0.015
R21878 VSS.n104 VSS.n103 0.015
R21879 VSS.n117 VSS.n115 0.015
R21880 VSS.n14093 VSS.n14092 0.015
R21881 VSS.n14094 VSS.n14093 0.015
R21882 VSS.n7073 VSS.n7072 0.015
R21883 VSS.n132 VSS.n130 0.015
R21884 VSS.n133 VSS.n132 0.015
R21885 VSS.n134 VSS.n133 0.015
R21886 VSS.n125 VSS.n124 0.015
R21887 VSS.n138 VSS.n136 0.015
R21888 VSS.n10575 VSS.n10574 0.015
R21889 VSS.n10576 VSS.n10575 0.015
R21890 VSS.n510 VSS.n509 0.015
R21891 VSS.n153 VSS.n151 0.015
R21892 VSS.n154 VSS.n153 0.015
R21893 VSS.n155 VSS.n154 0.015
R21894 VSS.n146 VSS.n145 0.015
R21895 VSS.n159 VSS.n157 0.015
R21896 VSS.n7056 VSS.n7055 0.015
R21897 VSS.n7057 VSS.n7056 0.015
R21898 VSS.n452 VSS.n451 0.015
R21899 VSS.n174 VSS.n172 0.015
R21900 VSS.n175 VSS.n174 0.015
R21901 VSS.n176 VSS.n175 0.015
R21902 VSS.n167 VSS.n166 0.015
R21903 VSS.n180 VSS.n178 0.015
R21904 VSS.n468 VSS.n467 0.015
R21905 VSS.n469 VSS.n468 0.015
R21906 VSS.n313 VSS.n312 0.015
R21907 VSS.n195 VSS.n193 0.015
R21908 VSS.n196 VSS.n195 0.015
R21909 VSS.n197 VSS.n196 0.015
R21910 VSS.n188 VSS.n187 0.015
R21911 VSS.n201 VSS.n199 0.015
R21912 VSS.n340 VSS.n339 0.015
R21913 VSS.n341 VSS.n340 0.015
R21914 VSS.n302 VSS.n301 0.015
R21915 VSS.n18256 VSS.n18254 0.015
R21916 VSS.n18235 VSS.n10 0.015
R21917 VSS.n18322 VSS.n18319 0.015
R21918 VSS.n496 VSS.n472 0.014
R21919 VSS.n18096 VSS.n18095 0.014
R21920 VSS.n17649 VSS.n17648 0.014
R21921 VSS.n17617 VSS.n17616 0.014
R21922 VSS.n14107 VSS.n14106 0.014
R21923 VSS.n10585 VSS.n10584 0.014
R21924 VSS.n7067 VSS.n7066 0.014
R21925 VSS.n504 VSS.n503 0.014
R21926 VSS.n446 VSS.n445 0.014
R21927 VSS.n17739 VSS.n17734 0.014
R21928 VSS.n18041 VSS.n18040 0.013
R21929 VSS.n18127 VSS.n18126 0.013
R21930 VSS.n269 VSS.n268 0.013
R21931 VSS.n220 VSS.n219 0.013
R21932 VSS.n18271 VSS.n18270 0.013
R21933 VSS.n5 VSS.n4 0.013
R21934 VSS.n22 VSS.n21 0.013
R21935 VSS.n48 VSS.n47 0.013
R21936 VSS.n17622 VSS.n17621 0.013
R21937 VSS.n67 VSS.n66 0.013
R21938 VSS.n14112 VSS.n14111 0.013
R21939 VSS.n88 VSS.n87 0.013
R21940 VSS.n10590 VSS.n10589 0.013
R21941 VSS.n109 VSS.n108 0.013
R21942 VSS.n7072 VSS.n7071 0.013
R21943 VSS.n130 VSS.n129 0.013
R21944 VSS.n509 VSS.n508 0.013
R21945 VSS.n151 VSS.n150 0.013
R21946 VSS.n451 VSS.n450 0.013
R21947 VSS.n172 VSS.n171 0.013
R21948 VSS.n312 VSS.n311 0.013
R21949 VSS.n193 VSS.n192 0.013
R21950 VSS.n301 VSS.n300 0.013
R21951 VSS.n18254 VSS.n18253 0.013
R21952 VSS.n10 VSS.n9 0.013
R21953 VSS.n18319 VSS.n18318 0.013
R21954 VSS.n251 VSS.n250 0.012
R21955 VSS.n253 VSS.n252 0.012
R21956 VSS.n18036 VSS.n18035 0.012
R21957 VSS.n18132 VSS.n18131 0.012
R21958 VSS.n18122 VSS.n18121 0.012
R21959 VSS.n14660 VSS.n14659 0.012
R21960 VSS.n14674 VSS.n14673 0.012
R21961 VSS.n14688 VSS.n14687 0.012
R21962 VSS.n14702 VSS.n14701 0.012
R21963 VSS.n14716 VSS.n14715 0.012
R21964 VSS.n14735 VSS.n14734 0.012
R21965 VSS.n14737 VSS.n14736 0.012
R21966 VSS.n14752 VSS.n14751 0.012
R21967 VSS.n14766 VSS.n14765 0.012
R21968 VSS.n14780 VSS.n14779 0.012
R21969 VSS.n14794 VSS.n14793 0.012
R21970 VSS.n14811 VSS.n14810 0.012
R21971 VSS.n14916 VSS.n14915 0.012
R21972 VSS.n14930 VSS.n14929 0.012
R21973 VSS.n14944 VSS.n14943 0.012
R21974 VSS.n14958 VSS.n14957 0.012
R21975 VSS.n14972 VSS.n14971 0.012
R21976 VSS.n14991 VSS.n14990 0.012
R21977 VSS.n14993 VSS.n14992 0.012
R21978 VSS.n15008 VSS.n15007 0.012
R21979 VSS.n15022 VSS.n15021 0.012
R21980 VSS.n15036 VSS.n15035 0.012
R21981 VSS.n15050 VSS.n15049 0.012
R21982 VSS.n15067 VSS.n15066 0.012
R21983 VSS.n15160 VSS.n15159 0.012
R21984 VSS.n15174 VSS.n15173 0.012
R21985 VSS.n15188 VSS.n15187 0.012
R21986 VSS.n15202 VSS.n15201 0.012
R21987 VSS.n15216 VSS.n15215 0.012
R21988 VSS.n15235 VSS.n15234 0.012
R21989 VSS.n15237 VSS.n15236 0.012
R21990 VSS.n15252 VSS.n15251 0.012
R21991 VSS.n15266 VSS.n15265 0.012
R21992 VSS.n15280 VSS.n15279 0.012
R21993 VSS.n15294 VSS.n15293 0.012
R21994 VSS.n15311 VSS.n15310 0.012
R21995 VSS.n15404 VSS.n15403 0.012
R21996 VSS.n15418 VSS.n15417 0.012
R21997 VSS.n15432 VSS.n15431 0.012
R21998 VSS.n15446 VSS.n15445 0.012
R21999 VSS.n15460 VSS.n15459 0.012
R22000 VSS.n15479 VSS.n15478 0.012
R22001 VSS.n15481 VSS.n15480 0.012
R22002 VSS.n15496 VSS.n15495 0.012
R22003 VSS.n15510 VSS.n15509 0.012
R22004 VSS.n15524 VSS.n15523 0.012
R22005 VSS.n15538 VSS.n15537 0.012
R22006 VSS.n15555 VSS.n15554 0.012
R22007 VSS.n15648 VSS.n15647 0.012
R22008 VSS.n15662 VSS.n15661 0.012
R22009 VSS.n15676 VSS.n15675 0.012
R22010 VSS.n15690 VSS.n15689 0.012
R22011 VSS.n15704 VSS.n15703 0.012
R22012 VSS.n15723 VSS.n15722 0.012
R22013 VSS.n15725 VSS.n15724 0.012
R22014 VSS.n15740 VSS.n15739 0.012
R22015 VSS.n15754 VSS.n15753 0.012
R22016 VSS.n15768 VSS.n15767 0.012
R22017 VSS.n15782 VSS.n15781 0.012
R22018 VSS.n15799 VSS.n15798 0.012
R22019 VSS.n15892 VSS.n15891 0.012
R22020 VSS.n15906 VSS.n15905 0.012
R22021 VSS.n15920 VSS.n15919 0.012
R22022 VSS.n15934 VSS.n15933 0.012
R22023 VSS.n15948 VSS.n15947 0.012
R22024 VSS.n15967 VSS.n15966 0.012
R22025 VSS.n15969 VSS.n15968 0.012
R22026 VSS.n15984 VSS.n15983 0.012
R22027 VSS.n15998 VSS.n15997 0.012
R22028 VSS.n16012 VSS.n16011 0.012
R22029 VSS.n16026 VSS.n16025 0.012
R22030 VSS.n16043 VSS.n16042 0.012
R22031 VSS.n16136 VSS.n16135 0.012
R22032 VSS.n16150 VSS.n16149 0.012
R22033 VSS.n16164 VSS.n16163 0.012
R22034 VSS.n16178 VSS.n16177 0.012
R22035 VSS.n16192 VSS.n16191 0.012
R22036 VSS.n16211 VSS.n16210 0.012
R22037 VSS.n16213 VSS.n16212 0.012
R22038 VSS.n16228 VSS.n16227 0.012
R22039 VSS.n16242 VSS.n16241 0.012
R22040 VSS.n16256 VSS.n16255 0.012
R22041 VSS.n16270 VSS.n16269 0.012
R22042 VSS.n16287 VSS.n16286 0.012
R22043 VSS.n16392 VSS.n16391 0.012
R22044 VSS.n16406 VSS.n16405 0.012
R22045 VSS.n16420 VSS.n16419 0.012
R22046 VSS.n16434 VSS.n16433 0.012
R22047 VSS.n16448 VSS.n16447 0.012
R22048 VSS.n16467 VSS.n16466 0.012
R22049 VSS.n16469 VSS.n16468 0.012
R22050 VSS.n16484 VSS.n16483 0.012
R22051 VSS.n16498 VSS.n16497 0.012
R22052 VSS.n16512 VSS.n16511 0.012
R22053 VSS.n16526 VSS.n16525 0.012
R22054 VSS.n16586 VSS.n16572 0.012
R22055 VSS.n14144 VSS.n14143 0.012
R22056 VSS.n14156 VSS.n14155 0.012
R22057 VSS.n14168 VSS.n14167 0.012
R22058 VSS.n14180 VSS.n14179 0.012
R22059 VSS.n14192 VSS.n14191 0.012
R22060 VSS.n14204 VSS.n14203 0.012
R22061 VSS.n14216 VSS.n14215 0.012
R22062 VSS.n14228 VSS.n14227 0.012
R22063 VSS.n14285 VSS.n14284 0.012
R22064 VSS.n14324 VSS.n14323 0.012
R22065 VSS.n14336 VSS.n14335 0.012
R22066 VSS.n14348 VSS.n14347 0.012
R22067 VSS.n14360 VSS.n14359 0.012
R22068 VSS.n14372 VSS.n14371 0.012
R22069 VSS.n14384 VSS.n14383 0.012
R22070 VSS.n14396 VSS.n14395 0.012
R22071 VSS.n14408 VSS.n14407 0.012
R22072 VSS.n14465 VSS.n14464 0.012
R22073 VSS.n17584 VSS.n17527 0.012
R22074 VSS.n17525 VSS.n17515 0.012
R22075 VSS.n17513 VSS.n17503 0.012
R22076 VSS.n17501 VSS.n17491 0.012
R22077 VSS.n17489 VSS.n17479 0.012
R22078 VSS.n17468 VSS.n17467 0.012
R22079 VSS.n17465 VSS.n17455 0.012
R22080 VSS.n17453 VSS.n17443 0.012
R22081 VSS.n17441 VSS.n17431 0.012
R22082 VSS.n17416 VSS.n17359 0.012
R22083 VSS.n17357 VSS.n17347 0.012
R22084 VSS.n17345 VSS.n17335 0.012
R22085 VSS.n17333 VSS.n17323 0.012
R22086 VSS.n17321 VSS.n17311 0.012
R22087 VSS.n17300 VSS.n17299 0.012
R22088 VSS.n17297 VSS.n17287 0.012
R22089 VSS.n17285 VSS.n17275 0.012
R22090 VSS.n17273 VSS.n17263 0.012
R22091 VSS.n17248 VSS.n17191 0.012
R22092 VSS.n17189 VSS.n17179 0.012
R22093 VSS.n17177 VSS.n17167 0.012
R22094 VSS.n17165 VSS.n17155 0.012
R22095 VSS.n17153 VSS.n17143 0.012
R22096 VSS.n17132 VSS.n17131 0.012
R22097 VSS.n17129 VSS.n17119 0.012
R22098 VSS.n17117 VSS.n17107 0.012
R22099 VSS.n17105 VSS.n17095 0.012
R22100 VSS.n17080 VSS.n17023 0.012
R22101 VSS.n17021 VSS.n17011 0.012
R22102 VSS.n17009 VSS.n16999 0.012
R22103 VSS.n16997 VSS.n16987 0.012
R22104 VSS.n16985 VSS.n16975 0.012
R22105 VSS.n16964 VSS.n16963 0.012
R22106 VSS.n16961 VSS.n16951 0.012
R22107 VSS.n16949 VSS.n16939 0.012
R22108 VSS.n16937 VSS.n16927 0.012
R22109 VSS.n16912 VSS.n16855 0.012
R22110 VSS.n16853 VSS.n16843 0.012
R22111 VSS.n16841 VSS.n16831 0.012
R22112 VSS.n16829 VSS.n16819 0.012
R22113 VSS.n16817 VSS.n16807 0.012
R22114 VSS.n16796 VSS.n16795 0.012
R22115 VSS.n16793 VSS.n16783 0.012
R22116 VSS.n16781 VSS.n16771 0.012
R22117 VSS.n16769 VSS.n16759 0.012
R22118 VSS.n16744 VSS.n16687 0.012
R22119 VSS.n16685 VSS.n16675 0.012
R22120 VSS.n16673 VSS.n16663 0.012
R22121 VSS.n16661 VSS.n16651 0.012
R22122 VSS.n16649 VSS.n16639 0.012
R22123 VSS.n16628 VSS.n16627 0.012
R22124 VSS.n16625 VSS.n16615 0.012
R22125 VSS.n16613 VSS.n16603 0.012
R22126 VSS.n16601 VSS.n16591 0.012
R22127 VSS.n16590 VSS.n16589 0.012
R22128 VSS.n10709 VSS.n10708 0.012
R22129 VSS.n10723 VSS.n10722 0.012
R22130 VSS.n10737 VSS.n10736 0.012
R22131 VSS.n10751 VSS.n10750 0.012
R22132 VSS.n10765 VSS.n10764 0.012
R22133 VSS.n10784 VSS.n10783 0.012
R22134 VSS.n10786 VSS.n10785 0.012
R22135 VSS.n10801 VSS.n10800 0.012
R22136 VSS.n10815 VSS.n10814 0.012
R22137 VSS.n10829 VSS.n10828 0.012
R22138 VSS.n10843 VSS.n10842 0.012
R22139 VSS.n10860 VSS.n10859 0.012
R22140 VSS.n10965 VSS.n10964 0.012
R22141 VSS.n10979 VSS.n10978 0.012
R22142 VSS.n10993 VSS.n10992 0.012
R22143 VSS.n11007 VSS.n11006 0.012
R22144 VSS.n11021 VSS.n11020 0.012
R22145 VSS.n11040 VSS.n11039 0.012
R22146 VSS.n11042 VSS.n11041 0.012
R22147 VSS.n11057 VSS.n11056 0.012
R22148 VSS.n11071 VSS.n11070 0.012
R22149 VSS.n11085 VSS.n11084 0.012
R22150 VSS.n11099 VSS.n11098 0.012
R22151 VSS.n11116 VSS.n11115 0.012
R22152 VSS.n11209 VSS.n11208 0.012
R22153 VSS.n11223 VSS.n11222 0.012
R22154 VSS.n11237 VSS.n11236 0.012
R22155 VSS.n11251 VSS.n11250 0.012
R22156 VSS.n11265 VSS.n11264 0.012
R22157 VSS.n11284 VSS.n11283 0.012
R22158 VSS.n11286 VSS.n11285 0.012
R22159 VSS.n11301 VSS.n11300 0.012
R22160 VSS.n11315 VSS.n11314 0.012
R22161 VSS.n11329 VSS.n11328 0.012
R22162 VSS.n11343 VSS.n11342 0.012
R22163 VSS.n11360 VSS.n11359 0.012
R22164 VSS.n11453 VSS.n11452 0.012
R22165 VSS.n11467 VSS.n11466 0.012
R22166 VSS.n11481 VSS.n11480 0.012
R22167 VSS.n11495 VSS.n11494 0.012
R22168 VSS.n11509 VSS.n11508 0.012
R22169 VSS.n11528 VSS.n11527 0.012
R22170 VSS.n11530 VSS.n11529 0.012
R22171 VSS.n11545 VSS.n11544 0.012
R22172 VSS.n11559 VSS.n11558 0.012
R22173 VSS.n11573 VSS.n11572 0.012
R22174 VSS.n11587 VSS.n11586 0.012
R22175 VSS.n11604 VSS.n11603 0.012
R22176 VSS.n11697 VSS.n11696 0.012
R22177 VSS.n11711 VSS.n11710 0.012
R22178 VSS.n11725 VSS.n11724 0.012
R22179 VSS.n11739 VSS.n11738 0.012
R22180 VSS.n11753 VSS.n11752 0.012
R22181 VSS.n11772 VSS.n11771 0.012
R22182 VSS.n11774 VSS.n11773 0.012
R22183 VSS.n11789 VSS.n11788 0.012
R22184 VSS.n11803 VSS.n11802 0.012
R22185 VSS.n11817 VSS.n11816 0.012
R22186 VSS.n11831 VSS.n11830 0.012
R22187 VSS.n11848 VSS.n11847 0.012
R22188 VSS.n11941 VSS.n11940 0.012
R22189 VSS.n11955 VSS.n11954 0.012
R22190 VSS.n11969 VSS.n11968 0.012
R22191 VSS.n11983 VSS.n11982 0.012
R22192 VSS.n11997 VSS.n11996 0.012
R22193 VSS.n12016 VSS.n12015 0.012
R22194 VSS.n12018 VSS.n12017 0.012
R22195 VSS.n12033 VSS.n12032 0.012
R22196 VSS.n12047 VSS.n12046 0.012
R22197 VSS.n12061 VSS.n12060 0.012
R22198 VSS.n12075 VSS.n12074 0.012
R22199 VSS.n12092 VSS.n12091 0.012
R22200 VSS.n12185 VSS.n12184 0.012
R22201 VSS.n12199 VSS.n12198 0.012
R22202 VSS.n12213 VSS.n12212 0.012
R22203 VSS.n12227 VSS.n12226 0.012
R22204 VSS.n12241 VSS.n12240 0.012
R22205 VSS.n12260 VSS.n12259 0.012
R22206 VSS.n12262 VSS.n12261 0.012
R22207 VSS.n12277 VSS.n12276 0.012
R22208 VSS.n12291 VSS.n12290 0.012
R22209 VSS.n12305 VSS.n12304 0.012
R22210 VSS.n12319 VSS.n12318 0.012
R22211 VSS.n12336 VSS.n12335 0.012
R22212 VSS.n12441 VSS.n12440 0.012
R22213 VSS.n12455 VSS.n12454 0.012
R22214 VSS.n12469 VSS.n12468 0.012
R22215 VSS.n12483 VSS.n12482 0.012
R22216 VSS.n12497 VSS.n12496 0.012
R22217 VSS.n12516 VSS.n12515 0.012
R22218 VSS.n12518 VSS.n12517 0.012
R22219 VSS.n12533 VSS.n12532 0.012
R22220 VSS.n12547 VSS.n12546 0.012
R22221 VSS.n12561 VSS.n12560 0.012
R22222 VSS.n12575 VSS.n12574 0.012
R22223 VSS.n12635 VSS.n12621 0.012
R22224 VSS.n12661 VSS.n12660 0.012
R22225 VSS.n12673 VSS.n12672 0.012
R22226 VSS.n12685 VSS.n12684 0.012
R22227 VSS.n12697 VSS.n12696 0.012
R22228 VSS.n12709 VSS.n12708 0.012
R22229 VSS.n12721 VSS.n12720 0.012
R22230 VSS.n12733 VSS.n12732 0.012
R22231 VSS.n12745 VSS.n12744 0.012
R22232 VSS.n12802 VSS.n12801 0.012
R22233 VSS.n12841 VSS.n12840 0.012
R22234 VSS.n12853 VSS.n12852 0.012
R22235 VSS.n12865 VSS.n12864 0.012
R22236 VSS.n12877 VSS.n12876 0.012
R22237 VSS.n12889 VSS.n12888 0.012
R22238 VSS.n12901 VSS.n12900 0.012
R22239 VSS.n12913 VSS.n12912 0.012
R22240 VSS.n12925 VSS.n12924 0.012
R22241 VSS.n12982 VSS.n12981 0.012
R22242 VSS.n13021 VSS.n13020 0.012
R22243 VSS.n13033 VSS.n13032 0.012
R22244 VSS.n13045 VSS.n13044 0.012
R22245 VSS.n13057 VSS.n13056 0.012
R22246 VSS.n13069 VSS.n13068 0.012
R22247 VSS.n13081 VSS.n13080 0.012
R22248 VSS.n13093 VSS.n13092 0.012
R22249 VSS.n13105 VSS.n13104 0.012
R22250 VSS.n13162 VSS.n13161 0.012
R22251 VSS.n13201 VSS.n13200 0.012
R22252 VSS.n13213 VSS.n13212 0.012
R22253 VSS.n13225 VSS.n13224 0.012
R22254 VSS.n13237 VSS.n13236 0.012
R22255 VSS.n13249 VSS.n13248 0.012
R22256 VSS.n13261 VSS.n13260 0.012
R22257 VSS.n13273 VSS.n13272 0.012
R22258 VSS.n13285 VSS.n13284 0.012
R22259 VSS.n13342 VSS.n13341 0.012
R22260 VSS.n13381 VSS.n13380 0.012
R22261 VSS.n13393 VSS.n13392 0.012
R22262 VSS.n13405 VSS.n13404 0.012
R22263 VSS.n13417 VSS.n13416 0.012
R22264 VSS.n13429 VSS.n13428 0.012
R22265 VSS.n13441 VSS.n13440 0.012
R22266 VSS.n13453 VSS.n13452 0.012
R22267 VSS.n13465 VSS.n13464 0.012
R22268 VSS.n13522 VSS.n13521 0.012
R22269 VSS.n13561 VSS.n13560 0.012
R22270 VSS.n13573 VSS.n13572 0.012
R22271 VSS.n13585 VSS.n13584 0.012
R22272 VSS.n13597 VSS.n13596 0.012
R22273 VSS.n13609 VSS.n13608 0.012
R22274 VSS.n13621 VSS.n13620 0.012
R22275 VSS.n13633 VSS.n13632 0.012
R22276 VSS.n13645 VSS.n13644 0.012
R22277 VSS.n13702 VSS.n13701 0.012
R22278 VSS.n13741 VSS.n13740 0.012
R22279 VSS.n13753 VSS.n13752 0.012
R22280 VSS.n13765 VSS.n13764 0.012
R22281 VSS.n13777 VSS.n13776 0.012
R22282 VSS.n13789 VSS.n13788 0.012
R22283 VSS.n13801 VSS.n13800 0.012
R22284 VSS.n13813 VSS.n13812 0.012
R22285 VSS.n13825 VSS.n13824 0.012
R22286 VSS.n13882 VSS.n13881 0.012
R22287 VSS.n13921 VSS.n13920 0.012
R22288 VSS.n13933 VSS.n13932 0.012
R22289 VSS.n13945 VSS.n13944 0.012
R22290 VSS.n13957 VSS.n13956 0.012
R22291 VSS.n13969 VSS.n13968 0.012
R22292 VSS.n13981 VSS.n13980 0.012
R22293 VSS.n13993 VSS.n13992 0.012
R22294 VSS.n14005 VSS.n14004 0.012
R22295 VSS.n14062 VSS.n14061 0.012
R22296 VSS.n7277 VSS.n7276 0.012
R22297 VSS.n7291 VSS.n7290 0.012
R22298 VSS.n7305 VSS.n7304 0.012
R22299 VSS.n7319 VSS.n7318 0.012
R22300 VSS.n7333 VSS.n7332 0.012
R22301 VSS.n7352 VSS.n7351 0.012
R22302 VSS.n7354 VSS.n7353 0.012
R22303 VSS.n7369 VSS.n7368 0.012
R22304 VSS.n7383 VSS.n7382 0.012
R22305 VSS.n7397 VSS.n7396 0.012
R22306 VSS.n7411 VSS.n7410 0.012
R22307 VSS.n7428 VSS.n7427 0.012
R22308 VSS.n7533 VSS.n7532 0.012
R22309 VSS.n7547 VSS.n7546 0.012
R22310 VSS.n7561 VSS.n7560 0.012
R22311 VSS.n7575 VSS.n7574 0.012
R22312 VSS.n7589 VSS.n7588 0.012
R22313 VSS.n7608 VSS.n7607 0.012
R22314 VSS.n7610 VSS.n7609 0.012
R22315 VSS.n7625 VSS.n7624 0.012
R22316 VSS.n7639 VSS.n7638 0.012
R22317 VSS.n7653 VSS.n7652 0.012
R22318 VSS.n7667 VSS.n7666 0.012
R22319 VSS.n7684 VSS.n7683 0.012
R22320 VSS.n7777 VSS.n7776 0.012
R22321 VSS.n7791 VSS.n7790 0.012
R22322 VSS.n7805 VSS.n7804 0.012
R22323 VSS.n7819 VSS.n7818 0.012
R22324 VSS.n7833 VSS.n7832 0.012
R22325 VSS.n7852 VSS.n7851 0.012
R22326 VSS.n7854 VSS.n7853 0.012
R22327 VSS.n7869 VSS.n7868 0.012
R22328 VSS.n7883 VSS.n7882 0.012
R22329 VSS.n7897 VSS.n7896 0.012
R22330 VSS.n7911 VSS.n7910 0.012
R22331 VSS.n7928 VSS.n7927 0.012
R22332 VSS.n8021 VSS.n8020 0.012
R22333 VSS.n8035 VSS.n8034 0.012
R22334 VSS.n8049 VSS.n8048 0.012
R22335 VSS.n8063 VSS.n8062 0.012
R22336 VSS.n8077 VSS.n8076 0.012
R22337 VSS.n8096 VSS.n8095 0.012
R22338 VSS.n8098 VSS.n8097 0.012
R22339 VSS.n8113 VSS.n8112 0.012
R22340 VSS.n8127 VSS.n8126 0.012
R22341 VSS.n8141 VSS.n8140 0.012
R22342 VSS.n8155 VSS.n8154 0.012
R22343 VSS.n8172 VSS.n8171 0.012
R22344 VSS.n8265 VSS.n8264 0.012
R22345 VSS.n8279 VSS.n8278 0.012
R22346 VSS.n8293 VSS.n8292 0.012
R22347 VSS.n8307 VSS.n8306 0.012
R22348 VSS.n8321 VSS.n8320 0.012
R22349 VSS.n8340 VSS.n8339 0.012
R22350 VSS.n8342 VSS.n8341 0.012
R22351 VSS.n8357 VSS.n8356 0.012
R22352 VSS.n8371 VSS.n8370 0.012
R22353 VSS.n8385 VSS.n8384 0.012
R22354 VSS.n8399 VSS.n8398 0.012
R22355 VSS.n8416 VSS.n8415 0.012
R22356 VSS.n8509 VSS.n8508 0.012
R22357 VSS.n8523 VSS.n8522 0.012
R22358 VSS.n8537 VSS.n8536 0.012
R22359 VSS.n8551 VSS.n8550 0.012
R22360 VSS.n8565 VSS.n8564 0.012
R22361 VSS.n8584 VSS.n8583 0.012
R22362 VSS.n8586 VSS.n8585 0.012
R22363 VSS.n8601 VSS.n8600 0.012
R22364 VSS.n8615 VSS.n8614 0.012
R22365 VSS.n8629 VSS.n8628 0.012
R22366 VSS.n8643 VSS.n8642 0.012
R22367 VSS.n8660 VSS.n8659 0.012
R22368 VSS.n8753 VSS.n8752 0.012
R22369 VSS.n8767 VSS.n8766 0.012
R22370 VSS.n8781 VSS.n8780 0.012
R22371 VSS.n8795 VSS.n8794 0.012
R22372 VSS.n8809 VSS.n8808 0.012
R22373 VSS.n8828 VSS.n8827 0.012
R22374 VSS.n8830 VSS.n8829 0.012
R22375 VSS.n8845 VSS.n8844 0.012
R22376 VSS.n8859 VSS.n8858 0.012
R22377 VSS.n8873 VSS.n8872 0.012
R22378 VSS.n8887 VSS.n8886 0.012
R22379 VSS.n8904 VSS.n8903 0.012
R22380 VSS.n9009 VSS.n9008 0.012
R22381 VSS.n9023 VSS.n9022 0.012
R22382 VSS.n9037 VSS.n9036 0.012
R22383 VSS.n9051 VSS.n9050 0.012
R22384 VSS.n9065 VSS.n9064 0.012
R22385 VSS.n9084 VSS.n9083 0.012
R22386 VSS.n9086 VSS.n9085 0.012
R22387 VSS.n9101 VSS.n9100 0.012
R22388 VSS.n9115 VSS.n9114 0.012
R22389 VSS.n9129 VSS.n9128 0.012
R22390 VSS.n9143 VSS.n9142 0.012
R22391 VSS.n9203 VSS.n9189 0.012
R22392 VSS.n10548 VSS.n10492 0.012
R22393 VSS.n10490 VSS.n10480 0.012
R22394 VSS.n10478 VSS.n10468 0.012
R22395 VSS.n10466 VSS.n10456 0.012
R22396 VSS.n10454 VSS.n10444 0.012
R22397 VSS.n10433 VSS.n10432 0.012
R22398 VSS.n10430 VSS.n10420 0.012
R22399 VSS.n10418 VSS.n10408 0.012
R22400 VSS.n10406 VSS.n10396 0.012
R22401 VSS.n10380 VSS.n10325 0.012
R22402 VSS.n10323 VSS.n10313 0.012
R22403 VSS.n10311 VSS.n10301 0.012
R22404 VSS.n10299 VSS.n10289 0.012
R22405 VSS.n10287 VSS.n10277 0.012
R22406 VSS.n10266 VSS.n10265 0.012
R22407 VSS.n10263 VSS.n10253 0.012
R22408 VSS.n10251 VSS.n10241 0.012
R22409 VSS.n10239 VSS.n10229 0.012
R22410 VSS.n10212 VSS.n10157 0.012
R22411 VSS.n10155 VSS.n10145 0.012
R22412 VSS.n10143 VSS.n10133 0.012
R22413 VSS.n10131 VSS.n10121 0.012
R22414 VSS.n10119 VSS.n10109 0.012
R22415 VSS.n10098 VSS.n10097 0.012
R22416 VSS.n10095 VSS.n10085 0.012
R22417 VSS.n10083 VSS.n10073 0.012
R22418 VSS.n10071 VSS.n10061 0.012
R22419 VSS.n10044 VSS.n9989 0.012
R22420 VSS.n9987 VSS.n9977 0.012
R22421 VSS.n9975 VSS.n9965 0.012
R22422 VSS.n9963 VSS.n9953 0.012
R22423 VSS.n9951 VSS.n9941 0.012
R22424 VSS.n9930 VSS.n9929 0.012
R22425 VSS.n9927 VSS.n9917 0.012
R22426 VSS.n9915 VSS.n9905 0.012
R22427 VSS.n9903 VSS.n9893 0.012
R22428 VSS.n9876 VSS.n9821 0.012
R22429 VSS.n9819 VSS.n9809 0.012
R22430 VSS.n9807 VSS.n9797 0.012
R22431 VSS.n9795 VSS.n9785 0.012
R22432 VSS.n9783 VSS.n9773 0.012
R22433 VSS.n9762 VSS.n9761 0.012
R22434 VSS.n9759 VSS.n9749 0.012
R22435 VSS.n9747 VSS.n9737 0.012
R22436 VSS.n9735 VSS.n9725 0.012
R22437 VSS.n9708 VSS.n9653 0.012
R22438 VSS.n9651 VSS.n9641 0.012
R22439 VSS.n9639 VSS.n9629 0.012
R22440 VSS.n9627 VSS.n9617 0.012
R22441 VSS.n9615 VSS.n9605 0.012
R22442 VSS.n9594 VSS.n9593 0.012
R22443 VSS.n9591 VSS.n9581 0.012
R22444 VSS.n9579 VSS.n9569 0.012
R22445 VSS.n9567 VSS.n9557 0.012
R22446 VSS.n9540 VSS.n9485 0.012
R22447 VSS.n9483 VSS.n9473 0.012
R22448 VSS.n9471 VSS.n9461 0.012
R22449 VSS.n9459 VSS.n9449 0.012
R22450 VSS.n9447 VSS.n9437 0.012
R22451 VSS.n9426 VSS.n9425 0.012
R22452 VSS.n9423 VSS.n9413 0.012
R22453 VSS.n9411 VSS.n9401 0.012
R22454 VSS.n9399 VSS.n9389 0.012
R22455 VSS.n9372 VSS.n9317 0.012
R22456 VSS.n9315 VSS.n9305 0.012
R22457 VSS.n9303 VSS.n9293 0.012
R22458 VSS.n9291 VSS.n9281 0.012
R22459 VSS.n9279 VSS.n9269 0.012
R22460 VSS.n9258 VSS.n9257 0.012
R22461 VSS.n9255 VSS.n9245 0.012
R22462 VSS.n9243 VSS.n9233 0.012
R22463 VSS.n9231 VSS.n9221 0.012
R22464 VSS.n9220 VSS.n9206 0.012
R22465 VSS.n3461 VSS.n3459 0.012
R22466 VSS.n3797 VSS.n3796 0.012
R22467 VSS.n3786 VSS.n3785 0.012
R22468 VSS.n3480 VSS.n3468 0.012
R22469 VSS.n3774 VSS.n3773 0.012
R22470 VSS.n3763 VSS.n3762 0.012
R22471 VSS.n3499 VSS.n3487 0.012
R22472 VSS.n3751 VSS.n3750 0.012
R22473 VSS.n3740 VSS.n3739 0.012
R22474 VSS.n3518 VSS.n3506 0.012
R22475 VSS.n3728 VSS.n3727 0.012
R22476 VSS.n3717 VSS.n3716 0.012
R22477 VSS.n3573 VSS.n3559 0.012
R22478 VSS.n3704 VSS.n3703 0.012
R22479 VSS.n3693 VSS.n3692 0.012
R22480 VSS.n3592 VSS.n3580 0.012
R22481 VSS.n3681 VSS.n3680 0.012
R22482 VSS.n3670 VSS.n3669 0.012
R22483 VSS.n3611 VSS.n3599 0.012
R22484 VSS.n3658 VSS.n3657 0.012
R22485 VSS.n3647 VSS.n3646 0.012
R22486 VSS.n3634 VSS.n3618 0.012
R22487 VSS.n3635 VSS.n3391 0.012
R22488 VSS.n3954 VSS.n3953 0.012
R22489 VSS.n3967 VSS.n3966 0.012
R22490 VSS.n3978 VSS.n3375 0.012
R22491 VSS.n3989 VSS.n3369 0.012
R22492 VSS.n3990 VSS.n3361 0.012
R22493 VSS.n4002 VSS.n4001 0.012
R22494 VSS.n4013 VSS.n3354 0.012
R22495 VSS.n4024 VSS.n3348 0.012
R22496 VSS.n4025 VSS.n3340 0.012
R22497 VSS.n4037 VSS.n4036 0.012
R22498 VSS.n4048 VSS.n3333 0.012
R22499 VSS.n4059 VSS.n3327 0.012
R22500 VSS.n4415 VSS.n4414 0.012
R22501 VSS.n4073 VSS.n4060 0.012
R22502 VSS.n4401 VSS.n4400 0.012
R22503 VSS.n4390 VSS.n4389 0.012
R22504 VSS.n4092 VSS.n4080 0.012
R22505 VSS.n4378 VSS.n4377 0.012
R22506 VSS.n4367 VSS.n4366 0.012
R22507 VSS.n4111 VSS.n4099 0.012
R22508 VSS.n4355 VSS.n4354 0.012
R22509 VSS.n4344 VSS.n4343 0.012
R22510 VSS.n4130 VSS.n4118 0.012
R22511 VSS.n4332 VSS.n4331 0.012
R22512 VSS.n4321 VSS.n4320 0.012
R22513 VSS.n4185 VSS.n4171 0.012
R22514 VSS.n4308 VSS.n4307 0.012
R22515 VSS.n4297 VSS.n4296 0.012
R22516 VSS.n4204 VSS.n4192 0.012
R22517 VSS.n4285 VSS.n4284 0.012
R22518 VSS.n4274 VSS.n4273 0.012
R22519 VSS.n4223 VSS.n4211 0.012
R22520 VSS.n4262 VSS.n4261 0.012
R22521 VSS.n4251 VSS.n4250 0.012
R22522 VSS.n4239 VSS.n4230 0.012
R22523 VSS.n4538 VSS.n3222 0.012
R22524 VSS.n4540 VSS.n3219 0.012
R22525 VSS.n4555 VSS.n3213 0.012
R22526 VSS.n4556 VSS.n3205 0.012
R22527 VSS.n4568 VSS.n4567 0.012
R22528 VSS.n4579 VSS.n3198 0.012
R22529 VSS.n4590 VSS.n3192 0.012
R22530 VSS.n4591 VSS.n3184 0.012
R22531 VSS.n4603 VSS.n4602 0.012
R22532 VSS.n4614 VSS.n3177 0.012
R22533 VSS.n4625 VSS.n3171 0.012
R22534 VSS.n4626 VSS.n3163 0.012
R22535 VSS.n4638 VSS.n4637 0.012
R22536 VSS.n4649 VSS.n4648 0.012
R22537 VSS.n4663 VSS.n4650 0.012
R22538 VSS.n5010 VSS.n5009 0.012
R22539 VSS.n4999 VSS.n4998 0.012
R22540 VSS.n4682 VSS.n4670 0.012
R22541 VSS.n4987 VSS.n4986 0.012
R22542 VSS.n4976 VSS.n4975 0.012
R22543 VSS.n4701 VSS.n4689 0.012
R22544 VSS.n4964 VSS.n4963 0.012
R22545 VSS.n4953 VSS.n4952 0.012
R22546 VSS.n4720 VSS.n4708 0.012
R22547 VSS.n4941 VSS.n4940 0.012
R22548 VSS.n4930 VSS.n4929 0.012
R22549 VSS.n4775 VSS.n4761 0.012
R22550 VSS.n4917 VSS.n4916 0.012
R22551 VSS.n4906 VSS.n4905 0.012
R22552 VSS.n4794 VSS.n4782 0.012
R22553 VSS.n4894 VSS.n4893 0.012
R22554 VSS.n4883 VSS.n4882 0.012
R22555 VSS.n4813 VSS.n4801 0.012
R22556 VSS.n4871 VSS.n4870 0.012
R22557 VSS.n4860 VSS.n4859 0.012
R22558 VSS.n4832 VSS.n4820 0.012
R22559 VSS.n4848 VSS.n4847 0.012
R22560 VSS.n4837 VSS.n3095 0.012
R22561 VSS.n2382 VSS.n2381 0.012
R22562 VSS.n2450 VSS.n2449 0.012
R22563 VSS.n2441 VSS.n2440 0.012
R22564 VSS.n2434 VSS.n2385 0.012
R22565 VSS.n2428 VSS.n2391 0.012
R22566 VSS.n2422 VSS.n2395 0.012
R22567 VSS.n2417 VSS.n2398 0.012
R22568 VSS.n2411 VSS.n2401 0.012
R22569 VSS.n2404 VSS.n2285 0.012
R22570 VSS.n2472 VSS.n2471 0.012
R22571 VSS.n2540 VSS.n2539 0.012
R22572 VSS.n2531 VSS.n2530 0.012
R22573 VSS.n2524 VSS.n2475 0.012
R22574 VSS.n2518 VSS.n2481 0.012
R22575 VSS.n2512 VSS.n2485 0.012
R22576 VSS.n2507 VSS.n2488 0.012
R22577 VSS.n2501 VSS.n2491 0.012
R22578 VSS.n2494 VSS.n2195 0.012
R22579 VSS.n2562 VSS.n2561 0.012
R22580 VSS.n2630 VSS.n2629 0.012
R22581 VSS.n2621 VSS.n2620 0.012
R22582 VSS.n2614 VSS.n2565 0.012
R22583 VSS.n2608 VSS.n2571 0.012
R22584 VSS.n2602 VSS.n2575 0.012
R22585 VSS.n2597 VSS.n2578 0.012
R22586 VSS.n2591 VSS.n2581 0.012
R22587 VSS.n2584 VSS.n2105 0.012
R22588 VSS.n2652 VSS.n2651 0.012
R22589 VSS.n2720 VSS.n2719 0.012
R22590 VSS.n2711 VSS.n2710 0.012
R22591 VSS.n2704 VSS.n2655 0.012
R22592 VSS.n2698 VSS.n2661 0.012
R22593 VSS.n2692 VSS.n2665 0.012
R22594 VSS.n2687 VSS.n2668 0.012
R22595 VSS.n2681 VSS.n2671 0.012
R22596 VSS.n2674 VSS.n2015 0.012
R22597 VSS.n2742 VSS.n2741 0.012
R22598 VSS.n2810 VSS.n2809 0.012
R22599 VSS.n2801 VSS.n2800 0.012
R22600 VSS.n2794 VSS.n2745 0.012
R22601 VSS.n2788 VSS.n2751 0.012
R22602 VSS.n2782 VSS.n2755 0.012
R22603 VSS.n2777 VSS.n2758 0.012
R22604 VSS.n2771 VSS.n2761 0.012
R22605 VSS.n2764 VSS.n1925 0.012
R22606 VSS.n2832 VSS.n2831 0.012
R22607 VSS.n2900 VSS.n2899 0.012
R22608 VSS.n2891 VSS.n2890 0.012
R22609 VSS.n2884 VSS.n2835 0.012
R22610 VSS.n2878 VSS.n2841 0.012
R22611 VSS.n2872 VSS.n2845 0.012
R22612 VSS.n2867 VSS.n2848 0.012
R22613 VSS.n2861 VSS.n2851 0.012
R22614 VSS.n2854 VSS.n1835 0.012
R22615 VSS.n2922 VSS.n2921 0.012
R22616 VSS.n2990 VSS.n2989 0.012
R22617 VSS.n2981 VSS.n2980 0.012
R22618 VSS.n2974 VSS.n2925 0.012
R22619 VSS.n2968 VSS.n2931 0.012
R22620 VSS.n2962 VSS.n2935 0.012
R22621 VSS.n2957 VSS.n2938 0.012
R22622 VSS.n2951 VSS.n2941 0.012
R22623 VSS.n2944 VSS.n1745 0.012
R22624 VSS.n3012 VSS.n3011 0.012
R22625 VSS.n3080 VSS.n3079 0.012
R22626 VSS.n3071 VSS.n3070 0.012
R22627 VSS.n3064 VSS.n3015 0.012
R22628 VSS.n3058 VSS.n3021 0.012
R22629 VSS.n3052 VSS.n3025 0.012
R22630 VSS.n3047 VSS.n3028 0.012
R22631 VSS.n3041 VSS.n3031 0.012
R22632 VSS.n3034 VSS.n1655 0.012
R22633 VSS.n5144 VSS.n1581 0.012
R22634 VSS.n5155 VSS.n1575 0.012
R22635 VSS.n5156 VSS.n1567 0.012
R22636 VSS.n5168 VSS.n5167 0.012
R22637 VSS.n5179 VSS.n1560 0.012
R22638 VSS.n5190 VSS.n1554 0.012
R22639 VSS.n5191 VSS.n1546 0.012
R22640 VSS.n5203 VSS.n5202 0.012
R22641 VSS.n5214 VSS.n1539 0.012
R22642 VSS.n5226 VSS.n1531 0.012
R22643 VSS.n5228 VSS.n1524 0.012
R22644 VSS.n5407 VSS.n5406 0.012
R22645 VSS.n5394 VSS.n5393 0.012
R22646 VSS.n5383 VSS.n5382 0.012
R22647 VSS.n5257 VSS.n5245 0.012
R22648 VSS.n5371 VSS.n5370 0.012
R22649 VSS.n5360 VSS.n5359 0.012
R22650 VSS.n5276 VSS.n5264 0.012
R22651 VSS.n5348 VSS.n5347 0.012
R22652 VSS.n5337 VSS.n5336 0.012
R22653 VSS.n5295 VSS.n5283 0.012
R22654 VSS.n5325 VSS.n5324 0.012
R22655 VSS.n5314 VSS.n5313 0.012
R22656 VSS.n5303 VSS.n5302 0.012
R22657 VSS.n5503 VSS.n1440 0.012
R22658 VSS.n5514 VSS.n1434 0.012
R22659 VSS.n5515 VSS.n1426 0.012
R22660 VSS.n5527 VSS.n5526 0.012
R22661 VSS.n5538 VSS.n1419 0.012
R22662 VSS.n5549 VSS.n1413 0.012
R22663 VSS.n5550 VSS.n1405 0.012
R22664 VSS.n5562 VSS.n5561 0.012
R22665 VSS.n5573 VSS.n1398 0.012
R22666 VSS.n5585 VSS.n1390 0.012
R22667 VSS.n5587 VSS.n1383 0.012
R22668 VSS.n5615 VSS.n5614 0.012
R22669 VSS.n5602 VSS.n519 0.012
R22670 VSS.n531 VSS.n520 0.012
R22671 VSS.n5773 VSS.n5772 0.012
R22672 VSS.n5762 VSS.n5761 0.012
R22673 VSS.n550 VSS.n538 0.012
R22674 VSS.n5750 VSS.n5749 0.012
R22675 VSS.n5739 VSS.n5738 0.012
R22676 VSS.n569 VSS.n557 0.012
R22677 VSS.n5727 VSS.n5726 0.012
R22678 VSS.n5716 VSS.n5715 0.012
R22679 VSS.n588 VSS.n576 0.012
R22680 VSS.n5704 VSS.n5703 0.012
R22681 VSS.n789 VSS.n777 0.012
R22682 VSS.n800 VSS.n771 0.012
R22683 VSS.n801 VSS.n763 0.012
R22684 VSS.n813 VSS.n812 0.012
R22685 VSS.n824 VSS.n756 0.012
R22686 VSS.n835 VSS.n750 0.012
R22687 VSS.n836 VSS.n742 0.012
R22688 VSS.n848 VSS.n847 0.012
R22689 VSS.n859 VSS.n735 0.012
R22690 VSS.n870 VSS.n729 0.012
R22691 VSS.n871 VSS.n720 0.012
R22692 VSS.n883 VSS.n882 0.012
R22693 VSS.n925 VSS.n924 0.012
R22694 VSS.n936 VSS.n705 0.012
R22695 VSS.n947 VSS.n699 0.012
R22696 VSS.n948 VSS.n691 0.012
R22697 VSS.n960 VSS.n959 0.012
R22698 VSS.n971 VSS.n684 0.012
R22699 VSS.n982 VSS.n678 0.012
R22700 VSS.n983 VSS.n670 0.012
R22701 VSS.n995 VSS.n994 0.012
R22702 VSS.n1006 VSS.n663 0.012
R22703 VSS.n1017 VSS.n657 0.012
R22704 VSS.n1264 VSS.n1263 0.012
R22705 VSS.n1031 VSS.n1018 0.012
R22706 VSS.n1250 VSS.n1249 0.012
R22707 VSS.n1239 VSS.n1238 0.012
R22708 VSS.n1050 VSS.n1038 0.012
R22709 VSS.n1227 VSS.n1226 0.012
R22710 VSS.n1216 VSS.n1215 0.012
R22711 VSS.n1069 VSS.n1057 0.012
R22712 VSS.n1204 VSS.n1203 0.012
R22713 VSS.n1193 VSS.n1192 0.012
R22714 VSS.n1088 VSS.n1076 0.012
R22715 VSS.n1181 VSS.n1180 0.012
R22716 VSS.n1170 VSS.n1169 0.012
R22717 VSS.n6676 VSS.n6675 0.012
R22718 VSS.n6743 VSS.n6742 0.012
R22719 VSS.n6734 VSS.n6733 0.012
R22720 VSS.n6727 VSS.n6679 0.012
R22721 VSS.n6721 VSS.n6685 0.012
R22722 VSS.n6715 VSS.n6689 0.012
R22723 VSS.n6709 VSS.n6693 0.012
R22724 VSS.n6704 VSS.n6696 0.012
R22725 VSS.n6699 VSS.n6579 0.012
R22726 VSS.n6766 VSS.n6765 0.012
R22727 VSS.n6833 VSS.n6832 0.012
R22728 VSS.n6824 VSS.n6823 0.012
R22729 VSS.n6817 VSS.n6769 0.012
R22730 VSS.n6811 VSS.n6775 0.012
R22731 VSS.n6805 VSS.n6779 0.012
R22732 VSS.n6799 VSS.n6783 0.012
R22733 VSS.n6794 VSS.n6786 0.012
R22734 VSS.n6789 VSS.n6489 0.012
R22735 VSS.n6856 VSS.n6855 0.012
R22736 VSS.n6923 VSS.n6922 0.012
R22737 VSS.n6914 VSS.n6913 0.012
R22738 VSS.n6907 VSS.n6859 0.012
R22739 VSS.n6901 VSS.n6865 0.012
R22740 VSS.n6895 VSS.n6869 0.012
R22741 VSS.n6889 VSS.n6873 0.012
R22742 VSS.n6884 VSS.n6876 0.012
R22743 VSS.n6879 VSS.n6399 0.012
R22744 VSS.n5793 VSS.n5786 0.012
R22745 VSS.n5799 VSS.n5798 0.012
R22746 VSS.n5805 VSS.n5804 0.012
R22747 VSS.n5811 VSS.n5810 0.012
R22748 VSS.n5816 VSS.n5815 0.012
R22749 VSS.n5823 VSS.n5822 0.012
R22750 VSS.n5829 VSS.n5828 0.012
R22751 VSS.n5835 VSS.n5834 0.012
R22752 VSS.n5840 VSS.n5839 0.012
R22753 VSS.n5900 VSS.n5893 0.012
R22754 VSS.n5908 VSS.n5891 0.012
R22755 VSS.n5916 VSS.n5889 0.012
R22756 VSS.n5924 VSS.n5887 0.012
R22757 VSS.n5932 VSS.n5885 0.012
R22758 VSS.n5940 VSS.n5883 0.012
R22759 VSS.n5948 VSS.n5881 0.012
R22760 VSS.n5956 VSS.n5879 0.012
R22761 VSS.n6371 VSS.n6370 0.012
R22762 VSS.n6016 VSS.n6009 0.012
R22763 VSS.n6024 VSS.n6007 0.012
R22764 VSS.n6032 VSS.n6005 0.012
R22765 VSS.n6040 VSS.n6003 0.012
R22766 VSS.n6048 VSS.n6001 0.012
R22767 VSS.n6056 VSS.n5999 0.012
R22768 VSS.n6064 VSS.n5997 0.012
R22769 VSS.n6072 VSS.n5995 0.012
R22770 VSS.n6307 VSS.n6306 0.012
R22771 VSS.n6132 VSS.n6125 0.012
R22772 VSS.n6140 VSS.n6123 0.012
R22773 VSS.n6148 VSS.n6121 0.012
R22774 VSS.n6156 VSS.n6119 0.012
R22775 VSS.n6164 VSS.n6117 0.012
R22776 VSS.n6172 VSS.n6115 0.012
R22777 VSS.n6180 VSS.n6113 0.012
R22778 VSS.n6188 VSS.n6111 0.012
R22779 VSS.n6243 VSS.n6242 0.012
R22780 VSS.n494 VSS.n472 0.012
R22781 VSS.n497 VSS.n496 0.011
R22782 VSS.n17765 VSS.n17743 0.011
R22783 VSS.n18095 VSS.n18094 0.01
R22784 VSS.n17648 VSS.n17647 0.01
R22785 VSS.n17616 VSS.n17615 0.01
R22786 VSS.n14106 VSS.n14105 0.01
R22787 VSS.n10584 VSS.n10583 0.01
R22788 VSS.n7066 VSS.n7065 0.01
R22789 VSS.n503 VSS.n502 0.01
R22790 VSS.n445 VSS.n444 0.01
R22791 VSS.n17739 VSS.n17738 0.01
R22792 VSS.n18032 VSS.n18031 0.01
R22793 VSS.n18132 VSS.n16 0.01
R22794 VSS.n18300 VSS.n18299 0.01
R22795 VSS.n18118 VSS.n18117 0.01
R22796 VSS.n14078 VSS.n14077 0.01
R22797 VSS.n7084 VSS.n7083 0.01
R22798 VSS.n398 VSS.n364 0.01
R22799 VSS.n417 VSS.n351 0.01
R22800 VSS.n18190 VSS.n18156 0.01
R22801 VSS.n18210 VSS.n18209 0.01
R22802 VSS.n18033 VSS.n18032 0.01
R22803 VSS.n18129 VSS.n18128 0.01
R22804 VSS.n18119 VSS.n18118 0.01
R22805 VSS.n18034 VSS.n18033 0.009
R22806 VSS.n18130 VSS.n18129 0.009
R22807 VSS.n18120 VSS.n18119 0.009
R22808 VSS.n273 VSS.n272 0.009
R22809 VSS.n265 VSS.n263 0.009
R22810 VSS.n278 VSS.n277 0.009
R22811 VSS.n289 VSS.n287 0.009
R22812 VSS.n274 VSS.n273 0.009
R22813 VSS.n287 VSS.n286 0.009
R22814 VSS.n226 VSS.n225 0.009
R22815 VSS.n215 VSS.n214 0.009
R22816 VSS.n229 VSS.n228 0.009
R22817 VSS.n213 VSS.n212 0.009
R22818 VSS.n232 VSS.n231 0.009
R22819 VSS.n210 VSS.n209 0.009
R22820 VSS.n239 VSS.n238 0.009
R22821 VSS.n222 VSS.n221 0.009
R22822 VSS.n341 VSS.n336 0.008
R22823 VSS.n469 VSS.n464 0.008
R22824 VSS.n7057 VSS.n7052 0.008
R22825 VSS.n10576 VSS.n10571 0.008
R22826 VSS.n14094 VSS.n14089 0.008
R22827 VSS.n17608 VSS.n17603 0.008
R22828 VSS.n17641 VSS.n17636 0.008
R22829 VSS.n18088 VSS.n36 0.008
R22830 VSS.n286 VSS.n284 0.008
R22831 VSS.n18100 VSS.n18099 0.008
R22832 VSS.n17655 VSS.n17654 0.008
R22833 VSS.n17666 VSS.n17665 0.008
R22834 VSS.n17676 VSS.n17675 0.008
R22835 VSS.n17687 VSS.n17686 0.008
R22836 VSS.n17698 VSS.n17697 0.008
R22837 VSS.n17709 VSS.n17708 0.008
R22838 VSS.n17719 VSS.n17718 0.008
R22839 VSS.n17730 VSS.n17729 0.008
R22840 VSS.n305 VSS.n304 0.008
R22841 VSS.n18039 VSS.n18038 0.008
R22842 VSS.n18037 VSS.n18036 0.008
R22843 VSS.n18125 VSS.n18124 0.008
R22844 VSS.n18123 VSS.n18122 0.008
R22845 VSS.n18303 VSS.n18302 0.008
R22846 VSS.n18305 VSS.n18304 0.008
R22847 VSS.n18308 VSS.n18307 0.008
R22848 VSS.n18310 VSS.n18309 0.008
R22849 VSS.n18313 VSS.n18312 0.008
R22850 VSS.n18315 VSS.n18314 0.008
R22851 VSS.n18323 VSS.n18322 0.008
R22852 VSS.n250 VSS.n249 0.008
R22853 VSS.n18236 VSS.n18235 0.008
R22854 VSS.n18238 VSS.n18237 0.008
R22855 VSS.n18241 VSS.n18240 0.008
R22856 VSS.n18243 VSS.n18242 0.008
R22857 VSS.n18246 VSS.n18245 0.008
R22858 VSS.n18248 VSS.n18247 0.008
R22859 VSS.n18257 VSS.n18250 0.008
R22860 VSS.n7046 VSS.n5785 0.008
R22861 VSS.n252 VSS.n251 0.007
R22862 VSS.n254 VSS.n253 0.007
R22863 VSS.n18035 VSS.n18034 0.007
R22864 VSS.n18121 VSS.n18120 0.007
R22865 VSS.n18131 VSS.n18130 0.007
R22866 VSS.n14098 VSS.n14097 0.006
R22867 VSS.n18096 VSS.n30 0.005
R22868 VSS.n18102 VSS.n18101 0.005
R22869 VSS.n29 VSS.n28 0.005
R22870 VSS.n26 VSS.n25 0.005
R22871 VSS.n18098 VSS.n18097 0.005
R22872 VSS.n24 VSS.n23 0.005
R22873 VSS.n17649 VSS.n17630 0.005
R22874 VSS.n17657 VSS.n17656 0.005
R22875 VSS.n17629 VSS.n17628 0.005
R22876 VSS.n17626 VSS.n17625 0.005
R22877 VSS.n17653 VSS.n17652 0.005
R22878 VSS.n17624 VSS.n17623 0.005
R22879 VSS.n17617 VSS.n14119 0.005
R22880 VSS.n17668 VSS.n17667 0.005
R22881 VSS.n14118 VSS.n14117 0.005
R22882 VSS.n14116 VSS.n14115 0.005
R22883 VSS.n17663 VSS.n17662 0.005
R22884 VSS.n14114 VSS.n14113 0.005
R22885 VSS.n14107 VSS.n10598 0.005
R22886 VSS.n17678 VSS.n17677 0.005
R22887 VSS.n10597 VSS.n10596 0.005
R22888 VSS.n10594 VSS.n10593 0.005
R22889 VSS.n17674 VSS.n17673 0.005
R22890 VSS.n10592 VSS.n10591 0.005
R22891 VSS.n10585 VSS.n7079 0.005
R22892 VSS.n17689 VSS.n17688 0.005
R22893 VSS.n7078 VSS.n7077 0.005
R22894 VSS.n7076 VSS.n7075 0.005
R22895 VSS.n17684 VSS.n17683 0.005
R22896 VSS.n7074 VSS.n7073 0.005
R22897 VSS.n7067 VSS.n516 0.005
R22898 VSS.n17700 VSS.n17699 0.005
R22899 VSS.n515 VSS.n514 0.005
R22900 VSS.n513 VSS.n512 0.005
R22901 VSS.n17695 VSS.n17694 0.005
R22902 VSS.n511 VSS.n510 0.005
R22903 VSS.n504 VSS.n458 0.005
R22904 VSS.n17711 VSS.n17710 0.005
R22905 VSS.n457 VSS.n456 0.005
R22906 VSS.n455 VSS.n454 0.005
R22907 VSS.n17706 VSS.n17705 0.005
R22908 VSS.n453 VSS.n452 0.005
R22909 VSS.n446 VSS.n320 0.005
R22910 VSS.n17721 VSS.n17720 0.005
R22911 VSS.n319 VSS.n318 0.005
R22912 VSS.n316 VSS.n315 0.005
R22913 VSS.n17717 VSS.n17716 0.005
R22914 VSS.n314 VSS.n313 0.005
R22915 VSS.n17734 VSS.n258 0.005
R22916 VSS.n17732 VSS.n17731 0.005
R22917 VSS.n307 VSS.n306 0.005
R22918 VSS.n17727 VSS.n17726 0.005
R22919 VSS.n303 VSS.n302 0.005
R22920 VSS.n400 VSS.n359 0.005
R22921 VSS.n410 VSS.n355 0.005
R22922 VSS.n18192 VSS.n18151 0.005
R22923 VSS.n18202 VSS.n18147 0.005
R22924 VSS.n14100 VSS.n14099 0.005
R22925 VSS.n247 VSS.n246 0.005
R22926 VSS.n3 VSS.n2 0.005
R22927 VSS.n34 VSS.n33 0.005
R22928 VSS.n17634 VSS.n17633 0.005
R22929 VSS.n17601 VSS.n17600 0.005
R22930 VSS.n14087 VSS.n14086 0.005
R22931 VSS.n10569 VSS.n10568 0.005
R22932 VSS.n7050 VSS.n7049 0.005
R22933 VSS.n462 VSS.n461 0.005
R22934 VSS.n334 VSS.n333 0.005
R22935 VSS.n234 VSS.n233 0.005
R22936 VSS.n18252 VSS.n18251 0.005
R22937 VSS.n14 VSS.n13 0.005
R22938 VSS.n18297 VSS.n18296 0.005
R22939 VSS.n10565 VSS.n10564 0.004
R22940 VSS.n238 VSS.n237 0.003
R22941 VSS.n272 VSS.n271 0.003
R22942 VSS.n18095 VSS.n18090 0.003
R22943 VSS.n18089 VSS.n18088 0.003
R22944 VSS.n17648 VSS.n17643 0.003
R22945 VSS.n17642 VSS.n17641 0.003
R22946 VSS.n17616 VSS.n17611 0.003
R22947 VSS.n17609 VSS.n17608 0.003
R22948 VSS.n14106 VSS.n14101 0.003
R22949 VSS.n14095 VSS.n14094 0.003
R22950 VSS.n10584 VSS.n10579 0.003
R22951 VSS.n10577 VSS.n10576 0.003
R22952 VSS.n7066 VSS.n7061 0.003
R22953 VSS.n7058 VSS.n7057 0.003
R22954 VSS.n503 VSS.n498 0.003
R22955 VSS.n470 VSS.n469 0.003
R22956 VSS.n445 VSS.n440 0.003
R22957 VSS.n342 VSS.n341 0.003
R22958 VSS.n17741 VSS.n17739 0.003
R22959 VSS.n18032 VSS.n18027 0.003
R22960 VSS.n18134 VSS.n18132 0.003
R22961 VSS.n18300 VSS.n18295 0.003
R22962 VSS.n18269 VSS.n18268 0.003
R22963 VSS.n267 VSS.n266 0.003
R22964 VSS.n18029 VSS.n18028 0.002
R22965 VSS.n18115 VSS.n18114 0.002
R22966 VSS.n20 VSS.n19 0.002
R22967 VSS.n17620 VSS.n17619 0.002
R22968 VSS.n14110 VSS.n14109 0.002
R22969 VSS.n10588 VSS.n10587 0.002
R22970 VSS.n7070 VSS.n7069 0.002
R22971 VSS.n507 VSS.n506 0.002
R22972 VSS.n449 VSS.n448 0.002
R22973 VSS.n310 VSS.n309 0.002
R22974 VSS.n299 VSS.n298 0.002
R22975 VSS.n46 VSS.n45 0.002
R22976 VSS.n65 VSS.n64 0.002
R22977 VSS.n86 VSS.n85 0.002
R22978 VSS.n107 VSS.n106 0.002
R22979 VSS.n128 VSS.n127 0.002
R22980 VSS.n149 VSS.n148 0.002
R22981 VSS.n170 VSS.n169 0.002
R22982 VSS.n191 VSS.n190 0.002
R22983 VSS.n218 VSS.n217 0.002
R22984 VSS.n18092 VSS.n18091 0.002
R22985 VSS.n17645 VSS.n17644 0.002
R22986 VSS.n17613 VSS.n17612 0.002
R22987 VSS.n14103 VSS.n14102 0.002
R22988 VSS.n10581 VSS.n10580 0.002
R22989 VSS.n7063 VSS.n7062 0.002
R22990 VSS.n500 VSS.n499 0.002
R22991 VSS.n442 VSS.n441 0.002
R22992 VSS.n17736 VSS.n17735 0.002
R22993 VSS.n17767 VSS.n17766 0.002
R22994 VSS.n18317 VSS.n18316 0.002
R22995 VSS.n282 VSS.n281 0.002
R22996 VSS.n8 VSS.n7 0.002
R22997 VSS.n242 VSS.n241 0.001
R22998 VSS.n18046 VSS.n18045 0.001
R22999 VSS.n18049 VSS.n18048 0.001
R23000 VSS.n18051 VSS.n18050 0.001
R23001 VSS.n18054 VSS.n18053 0.001
R23002 VSS.n18056 VSS.n18055 0.001
R23003 VSS.n18059 VSS.n18058 0.001
R23004 VSS.n18061 VSS.n18060 0.001
R23005 VSS.n18064 VSS.n18063 0.001
R23006 VSS.n18066 VSS.n18065 0.001
R23007 VSS.n18069 VSS.n18068 0.001
R23008 VSS.n18071 VSS.n18070 0.001
R23009 VSS.n18074 VSS.n18073 0.001
R23010 VSS.n18076 VSS.n18075 0.001
R23011 VSS.n18079 VSS.n18078 0.001
R23012 VSS.n18081 VSS.n18080 0.001
R23013 VSS.n40 VSS.n39 0.001
R23014 VSS.n18260 VSS.n18259 0.001
R23015 VSS.n18262 VSS.n18261 0.001
R23016 VSS.n18044 VSS.n18043 0.001
R23017 VSS.n38 VSS.n6 0.001
R23018 VSS.n294 VSS.n293 0.001
R23019 VSS.n18109 VSS.n18108 0.001
R23020 VSS.n18326 VSS.n18325 0.001
R23021 VSS.n268 VSS.n267 0.001
R23022 VSS.n283 VSS.n282 0.001
R23023 VSS.n219 VSS.n218 0.001
R23024 VSS.n235 VSS.n234 0.001
R23025 VSS.n18270 VSS.n18269 0.001
R23026 VSS.n4 VSS.n3 0.001
R23027 VSS.n18093 VSS.n18092 0.001
R23028 VSS.n21 VSS.n20 0.001
R23029 VSS.n47 VSS.n46 0.001
R23030 VSS.n35 VSS.n34 0.001
R23031 VSS.n17646 VSS.n17645 0.001
R23032 VSS.n17621 VSS.n17620 0.001
R23033 VSS.n66 VSS.n65 0.001
R23034 VSS.n17635 VSS.n17634 0.001
R23035 VSS.n17614 VSS.n17613 0.001
R23036 VSS.n14111 VSS.n14110 0.001
R23037 VSS.n87 VSS.n86 0.001
R23038 VSS.n17602 VSS.n17601 0.001
R23039 VSS.n14081 VSS.n14078 0.001
R23040 VSS.n14104 VSS.n14103 0.001
R23041 VSS.n10589 VSS.n10588 0.001
R23042 VSS.n108 VSS.n107 0.001
R23043 VSS.n14088 VSS.n14087 0.001
R23044 VSS.n10582 VSS.n10581 0.001
R23045 VSS.n7071 VSS.n7070 0.001
R23046 VSS.n129 VSS.n128 0.001
R23047 VSS.n10570 VSS.n10569 0.001
R23048 VSS.n7064 VSS.n7063 0.001
R23049 VSS.n508 VSS.n507 0.001
R23050 VSS.n150 VSS.n149 0.001
R23051 VSS.n7051 VSS.n7050 0.001
R23052 VSS.n501 VSS.n500 0.001
R23053 VSS.n450 VSS.n449 0.001
R23054 VSS.n171 VSS.n170 0.001
R23055 VSS.n463 VSS.n462 0.001
R23056 VSS.n443 VSS.n442 0.001
R23057 VSS.n311 VSS.n310 0.001
R23058 VSS.n192 VSS.n191 0.001
R23059 VSS.n335 VSS.n334 0.001
R23060 VSS.n17737 VSS.n17736 0.001
R23061 VSS.n300 VSS.n299 0.001
R23062 VSS.n248 VSS.n247 0.001
R23063 VSS.n18030 VSS.n18029 0.001
R23064 VSS.n240 VSS.n207 0.001
R23065 VSS.n18253 VSS.n18252 0.001
R23066 VSS.n9 VSS.n8 0.001
R23067 VSS.n15 VSS.n14 0.001
R23068 VSS.n18116 VSS.n18115 0.001
R23069 VSS.n18298 VSS.n18297 0.001
R23070 VSS.n18318 VSS.n18317 0.001
R23071 VSS.n17733 VSS.n17725 0.001
R23072 VSS.n17722 VSS.n17715 0.001
R23073 VSS.n17712 VSS.n17704 0.001
R23074 VSS.n17701 VSS.n17693 0.001
R23075 VSS.n17690 VSS.n17682 0.001
R23076 VSS.n17679 VSS.n17672 0.001
R23077 VSS.n17669 VSS.n17661 0.001
R23078 VSS.n17658 VSS.n17651 0.001
R23079 VSS.n18104 VSS.n18103 0.001
R23080 VSS.n18042 VSS.n244 0.001
R23081 VSS.n18264 VSS.n18263 0.001
R23082 VSS.n244 VSS.n243 0.001
R23083 VSS.n18285 VSS.n18264 0.001
R23084 VSS.n292 VSS.n262 0.001
R23085 VSS.n17733 VSS.n296 0.001
R23086 VSS.n17723 VSS.n17722 0.001
R23087 VSS.n17713 VSS.n17712 0.001
R23088 VSS.n17702 VSS.n17701 0.001
R23089 VSS.n17691 VSS.n17690 0.001
R23090 VSS.n17680 VSS.n17679 0.001
R23091 VSS.n17670 VSS.n17669 0.001
R23092 VSS.n17659 VSS.n17658 0.001
R23093 VSS.n18103 VSS.n17 0.001
R23094 VSS.n18110 VSS.n18106 0.001
R23095 VSS.n18324 VSS.n1 0.001
R23096 VSS.n18107 VSS.n1 0.001
R23097 VSS.n18106 VSS.n18105 0.001
R23098 VSS.n17650 VSS.n17 0.001
R23099 VSS.n17660 VSS.n17659 0.001
R23100 VSS.n17671 VSS.n17670 0.001
R23101 VSS.n17681 VSS.n17680 0.001
R23102 VSS.n17692 VSS.n17691 0.001
R23103 VSS.n17703 VSS.n17702 0.001
R23104 VSS.n17714 VSS.n17713 0.001
R23105 VSS.n17724 VSS.n17723 0.001
R23106 VSS.n296 VSS.n295 0.001
R23107 VSS.n262 VSS.n261 0.001
R23108 VSS.n18043 VSS.n18042 0.001
R23109 VSS.n18258 VSS.n6 0.001
R23110 VSS.n18047 VSS.n18046 0.001
R23111 VSS.n18048 VSS.n18047 0.001
R23112 VSS.n18052 VSS.n18051 0.001
R23113 VSS.n18053 VSS.n18052 0.001
R23114 VSS.n18057 VSS.n18056 0.001
R23115 VSS.n18058 VSS.n18057 0.001
R23116 VSS.n18062 VSS.n18061 0.001
R23117 VSS.n18063 VSS.n18062 0.001
R23118 VSS.n18067 VSS.n18066 0.001
R23119 VSS.n18068 VSS.n18067 0.001
R23120 VSS.n18072 VSS.n18071 0.001
R23121 VSS.n18073 VSS.n18072 0.001
R23122 VSS.n18077 VSS.n18076 0.001
R23123 VSS.n18078 VSS.n18077 0.001
R23124 VSS.n18082 VSS.n18081 0.001
R23125 VSS.n18082 VSS.n40 0.001
R23126 VSS.n18285 VSS.n18262 0.001
R23127 VSS.n241 VSS.n240 0.001
R23128 VSS.n18259 VSS.n18258 0.001
R23129 VSS.n18325 VSS.n18324 0.001
R23130 VSS.n18110 VSS.n18109 0.001
R23131 VSS.n293 VSS.n292 0.001
R23132 VSS.n18250 VSS.n18249 0.001
R23133 VSS.n18240 VSS.n18239 0.001
R23134 VSS.n228 VSS.n227 0.001
R23135 VSS.n212 VSS.n211 0.001
R23136 VSS.n18267 VSS.n18266 0.001
R23137 VSS.n18282 VSS.n18281 0.001
R23138 VSS.n58 VSS.n57 0.001
R23139 VSS.n56 VSS.n55 0.001
R23140 VSS.n77 VSS.n76 0.001
R23141 VSS.n75 VSS.n74 0.001
R23142 VSS.n98 VSS.n97 0.001
R23143 VSS.n96 VSS.n95 0.001
R23144 VSS.n119 VSS.n118 0.001
R23145 VSS.n117 VSS.n116 0.001
R23146 VSS.n140 VSS.n139 0.001
R23147 VSS.n138 VSS.n137 0.001
R23148 VSS.n161 VSS.n160 0.001
R23149 VSS.n159 VSS.n158 0.001
R23150 VSS.n182 VSS.n181 0.001
R23151 VSS.n180 VSS.n179 0.001
R23152 VSS.n203 VSS.n202 0.001
R23153 VSS.n201 VSS.n200 0.001
R23154 VSS.n17729 VSS.n17728 0.001
R23155 VSS.n18038 VSS.n256 0.001
R23156 VSS.n18040 VSS.n255 0.001
R23157 VSS.n18126 VSS.n18111 0.001
R23158 VSS.n18124 VSS.n18112 0.001
R23159 VSS.n18302 VSS.n18301 0.001
R23160 VSS.n18312 VSS.n18311 0.001
R23161 VSS.n18245 VSS.n18244 0.001
R23162 VSS.n18307 VSS.n18306 0.001
R23163 VSS.n18277 VSS.n18276 0.001
R23164 VSS.n18322 VSS.n18321 0.001
R23165 VSS.n14458 VSS.n14457 0.001
R23166 VSS.n14457 VSS.t10 0.001
R23167 VSS.n14278 VSS.n14277 0.001
R23168 VSS.n14277 VSS.t8 0.001
R23169 VSS.n14055 VSS.n14054 0.001
R23170 VSS.n14054 VSS.t32 0.001
R23171 VSS.n13875 VSS.n13874 0.001
R23172 VSS.n13874 VSS.t46 0.001
R23173 VSS.n13695 VSS.n13694 0.001
R23174 VSS.n13694 VSS.t44 0.001
R23175 VSS.n13515 VSS.n13514 0.001
R23176 VSS.n13514 VSS.t36 0.001
R23177 VSS.n13335 VSS.n13334 0.001
R23178 VSS.n13334 VSS.t34 0.001
R23179 VSS.n13155 VSS.n13154 0.001
R23180 VSS.n13154 VSS.t38 0.001
R23181 VSS.n12975 VSS.n12974 0.001
R23182 VSS.n12974 VSS.t42 0.001
R23183 VSS.n12795 VSS.n12794 0.001
R23184 VSS.n12794 VSS.t40 0.001
R23185 VSS.n9366 VSS.n9365 0.001
R23186 VSS.n9365 VSS.t48 0.001
R23187 VSS.n9534 VSS.n9533 0.001
R23188 VSS.n9533 VSS.t62 0.001
R23189 VSS.n9702 VSS.n9701 0.001
R23190 VSS.n9701 VSS.t60 0.001
R23191 VSS.n9870 VSS.n9869 0.001
R23192 VSS.n9869 VSS.t52 0.001
R23193 VSS.n10038 VSS.n10037 0.001
R23194 VSS.n10037 VSS.t50 0.001
R23195 VSS.n10206 VSS.n10205 0.001
R23196 VSS.n10205 VSS.t54 0.001
R23197 VSS.n10374 VSS.n10373 0.001
R23198 VSS.n10373 VSS.t58 0.001
R23199 VSS.n2458 VSS.n2307 0.001
R23200 VSS.t24 VSS.n2307 0.001
R23201 VSS.n2548 VSS.n2217 0.001
R23202 VSS.t26 VSS.n2217 0.001
R23203 VSS.n2638 VSS.n2127 0.001
R23204 VSS.t22 VSS.n2127 0.001
R23205 VSS.n2728 VSS.n2037 0.001
R23206 VSS.t18 VSS.n2037 0.001
R23207 VSS.n2818 VSS.n1947 0.001
R23208 VSS.t20 VSS.n1947 0.001
R23209 VSS.n2908 VSS.n1857 0.001
R23210 VSS.t28 VSS.n1857 0.001
R23211 VSS.n2998 VSS.n1767 0.001
R23212 VSS.t30 VSS.n1767 0.001
R23213 VSS.n3088 VSS.n1677 0.001
R23214 VSS.t16 VSS.n1677 0.001
R23215 VSS.n6932 VSS.n6421 0.001
R23216 VSS.t66 VSS.n6421 0.001
R23217 VSS.n6842 VSS.n6511 0.001
R23218 VSS.t70 VSS.n6511 0.001
R23219 VSS.n6752 VSS.n6601 0.001
R23220 VSS.t72 VSS.n6601 0.001
R23221 VSS.n18235 VSS.n18234 0.001
R23222 VSS.n18291 VSS.n18290 0.001
R23223 vbg.n172 vbg.n171 1412.31
R23224 vbg.n95 vbg.n92 176.62
R23225 vbg.n172 vbg 92.08
R23226 vbg.n0 vbg 60.003
R23227 vbg.n78 vbg.n77 54.344
R23228 vbg.n95 vbg.n94 54.344
R23229 vbg.n67 vbg.n66 47.551
R23230 vbg.n106 vbg.n105 47.551
R23231 vbg.n11 vbg.n10 44.155
R23232 vbg.n160 vbg.n159 44.155
R23233 vbg.n56 vbg.n55 40.758
R23234 vbg.n117 vbg.n116 40.758
R23235 vbg.n22 vbg.n21 37.362
R23236 vbg.n149 vbg.n148 37.362
R23237 vbg.n45 vbg.n44 33.965
R23238 vbg.n128 vbg.n127 33.965
R23239 vbg.n33 vbg.n32 30.568
R23240 vbg.n138 vbg.n137 30.568
R23241 vbg.n34 vbg.n33 27.172
R23242 vbg.n139 vbg.n138 27.172
R23243 vbg.n44 vbg.n43 23.775
R23244 vbg.n127 vbg.n126 23.775
R23245 vbg.n23 vbg.n22 20.379
R23246 vbg.n150 vbg.n149 20.379
R23247 vbg.n55 vbg.n54 16.982
R23248 vbg.n116 vbg.n115 16.982
R23249 vbg.n12 vbg.n11 13.586
R23250 vbg.n161 vbg.n160 13.586
R23251 vbg.n86 vbg.n85 13.176
R23252 vbg.n66 vbg.n65 10.189
R23253 vbg.n105 vbg.n104 10.189
R23254 vbg.n167 vbg.n166 9.3
R23255 vbg.n156 vbg.n155 9.3
R23256 vbg.n145 vbg.n144 9.3
R23257 vbg.n134 vbg.n133 9.3
R23258 vbg.n123 vbg.n122 9.3
R23259 vbg.n112 vbg.n111 9.3
R23260 vbg.n101 vbg.n100 9.3
R23261 vbg.n89 vbg.n88 9.3
R23262 vbg.n82 vbg.n81 9.3
R23263 vbg.n71 vbg.n70 9.3
R23264 vbg.n60 vbg.n59 9.3
R23265 vbg.n49 vbg.n48 9.3
R23266 vbg.n38 vbg.n37 9.3
R23267 vbg.n27 vbg.n26 9.3
R23268 vbg.n16 vbg.n15 9.3
R23269 vbg.n3 vbg.n2 9.3
R23270 vbg.n170 vbg.n169 9.3
R23271 vbg.n165 vbg.n164 9.3
R23272 vbg.n163 vbg.n162 9.3
R23273 vbg.n162 vbg.n161 9.3
R23274 vbg.n154 vbg.n153 9.3
R23275 vbg.n152 vbg.n151 9.3
R23276 vbg.n151 vbg.n150 9.3
R23277 vbg.n143 vbg.n142 9.3
R23278 vbg.n141 vbg.n140 9.3
R23279 vbg.n140 vbg.n139 9.3
R23280 vbg.n132 vbg.n131 9.3
R23281 vbg.n130 vbg.n129 9.3
R23282 vbg.n129 vbg.n128 9.3
R23283 vbg.n121 vbg.n120 9.3
R23284 vbg.n119 vbg.n118 9.3
R23285 vbg.n118 vbg.n117 9.3
R23286 vbg.n110 vbg.n109 9.3
R23287 vbg.n108 vbg.n107 9.3
R23288 vbg.n107 vbg.n106 9.3
R23289 vbg.n99 vbg.n98 9.3
R23290 vbg.n97 vbg.n96 9.3
R23291 vbg.n96 vbg.n95 9.3
R23292 vbg.n87 vbg.n86 9.3
R23293 vbg.n84 vbg.n83 9.3
R23294 vbg.n80 vbg.n79 9.3
R23295 vbg.n79 vbg.n78 9.3
R23296 vbg.n73 vbg.n72 9.3
R23297 vbg.n69 vbg.n68 9.3
R23298 vbg.n68 vbg.n67 9.3
R23299 vbg.n62 vbg.n61 9.3
R23300 vbg.n58 vbg.n57 9.3
R23301 vbg.n57 vbg.n56 9.3
R23302 vbg.n51 vbg.n50 9.3
R23303 vbg.n47 vbg.n46 9.3
R23304 vbg.n46 vbg.n45 9.3
R23305 vbg.n40 vbg.n39 9.3
R23306 vbg.n36 vbg.n35 9.3
R23307 vbg.n35 vbg.n34 9.3
R23308 vbg.n29 vbg.n28 9.3
R23309 vbg.n25 vbg.n24 9.3
R23310 vbg.n24 vbg.n23 9.3
R23311 vbg.n18 vbg.n17 9.3
R23312 vbg.n14 vbg.n13 9.3
R23313 vbg.n13 vbg.n12 9.3
R23314 vbg.n7 vbg.n6 9.3
R23315 vbg.n5 vbg.n4 9.3
R23316 vbg.n79 vbg.n75 6.023
R23317 vbg.n96 vbg.n91 6.023
R23318 vbg.n68 vbg.n64 5.27
R23319 vbg.n107 vbg.n103 5.27
R23320 vbg.n9 vbg.n8 4.894
R23321 vbg.n158 vbg.n157 4.894
R23322 vbg.n171 vbg.n170 4.84
R23323 vbg.n57 vbg.n53 4.517
R23324 vbg.n118 vbg.n114 4.517
R23325 vbg.n20 vbg.n19 4.141
R23326 vbg.n147 vbg.n146 4.141
R23327 vbg.n46 vbg.n42 3.764
R23328 vbg.n129 vbg.n125 3.764
R23329 vbg.n77 vbg.n76 3.396
R23330 vbg.n94 vbg.n93 3.396
R23331 vbg.n31 vbg.n30 3.388
R23332 vbg.n136 vbg.n135 3.388
R23333 vbg.n35 vbg.n31 3.011
R23334 vbg.n140 vbg.n136 3.011
R23335 vbg.n42 vbg.n41 2.635
R23336 vbg.n125 vbg.n124 2.635
R23337 vbg.n24 vbg.n20 2.258
R23338 vbg.n151 vbg.n147 2.258
R23339 vbg.n53 vbg.n52 1.882
R23340 vbg.n114 vbg.n113 1.882
R23341 vbg.n13 vbg.n9 1.505
R23342 vbg.n162 vbg.n158 1.505
R23343 vbg.n64 vbg.n63 1.129
R23344 vbg.n103 vbg.n102 1.129
R23345 vbg vbg.n172 0.853
R23346 vbg.n2 vbg.n1 0.851
R23347 vbg.n169 vbg.n168 0.851
R23348 vbg.n75 vbg.n74 0.376
R23349 vbg.n91 vbg.n90 0.376
R23350 vbg.n87 vbg.n84 0.19
R23351 vbg.n3 vbg.n0 0.152
R23352 vbg.n14 vbg.n7 0.144
R23353 vbg.n25 vbg.n18 0.144
R23354 vbg.n36 vbg.n29 0.144
R23355 vbg.n47 vbg.n40 0.144
R23356 vbg.n58 vbg.n51 0.144
R23357 vbg.n69 vbg.n62 0.144
R23358 vbg.n80 vbg.n73 0.144
R23359 vbg.n99 vbg.n97 0.144
R23360 vbg.n110 vbg.n108 0.144
R23361 vbg.n121 vbg.n119 0.144
R23362 vbg.n132 vbg.n130 0.144
R23363 vbg.n143 vbg.n141 0.144
R23364 vbg.n154 vbg.n152 0.144
R23365 vbg.n165 vbg.n163 0.144
R23366 vbg.n82 vbg.n80 0.043
R23367 vbg.n97 vbg.n89 0.043
R23368 vbg.n7 vbg.n5 0.04
R23369 vbg.n167 vbg.n165 0.04
R23370 vbg.n71 vbg.n69 0.038
R23371 vbg.n108 vbg.n101 0.038
R23372 vbg.n18 vbg.n16 0.035
R23373 vbg.n156 vbg.n154 0.035
R23374 vbg.n60 vbg.n58 0.032
R23375 vbg.n119 vbg.n112 0.032
R23376 vbg.n29 vbg.n27 0.029
R23377 vbg.n145 vbg.n143 0.029
R23378 vbg.n49 vbg.n47 0.027
R23379 vbg.n130 vbg.n123 0.027
R23380 vbg.n40 vbg.n38 0.024
R23381 vbg.n134 vbg.n132 0.024
R23382 vbg.n38 vbg.n36 0.021
R23383 vbg.n141 vbg.n134 0.021
R23384 vbg.n51 vbg.n49 0.019
R23385 vbg.n123 vbg.n121 0.019
R23386 vbg.n27 vbg.n25 0.016
R23387 vbg.n152 vbg.n145 0.016
R23388 vbg.n62 vbg.n60 0.013
R23389 vbg.n112 vbg.n110 0.013
R23390 vbg.n16 vbg.n14 0.01
R23391 vbg.n163 vbg.n156 0.01
R23392 vbg.n73 vbg.n71 0.008
R23393 vbg.n101 vbg.n99 0.008
R23394 vbg.n5 vbg.n3 0.005
R23395 vbg.n170 vbg.n167 0.005
R23396 vbg.n84 vbg.n82 0.002
R23397 vbg.n89 vbg.n87 0.002
R23398 VDD.n832 VDD 7803.62
R23399 VDD.n1506 VDD 7803.18
R23400 VDD.n443 VDD 7182.72
R23401 VDD.n188 VDD.n187 6898.54
R23402 VDD.n191 VDD.n189 6898.54
R23403 VDD.n902 VDD.n901 6713.54
R23404 VDD.n845 VDD.n844 6713.54
R23405 VDD.n643 VDD.t34 6271.13
R23406 VDD.n868 VDD 1647.66
R23407 VDD.n443 VDD.n442 1494.96
R23408 VDD.n1525 VDD 1077.32
R23409 VDD.n902 VDD 1077.32
R23410 VDD.n845 VDD 1077.32
R23411 VDD.n643 VDD 1077.32
R23412 VDD.n622 VDD 1077.32
R23413 VDD.n188 VDD 1077.32
R23414 VDD.n191 VDD 1077.32
R23415 VDD.n886 VDD.n870 934.848
R23416 VDD.n715 VDD.n714 934.848
R23417 VDD.n901 VDD.n870 749.848
R23418 VDD.n714 VDD.n713 749.848
R23419 VDD.n713 VDD.n703 749.848
R23420 VDD.n753 VDD.n703 749.848
R23421 VDD.n754 VDD.n753 749.848
R23422 VDD.n754 VDD.n696 749.848
R23423 VDD.n772 VDD.n696 749.848
R23424 VDD.n773 VDD.n772 749.848
R23425 VDD.n773 VDD.n690 749.848
R23426 VDD.n788 VDD.n690 749.848
R23427 VDD.n792 VDD.n788 749.848
R23428 VDD.n792 VDD.n791 749.848
R23429 VDD.n791 VDD.n790 749.848
R23430 VDD.n790 VDD.n789 749.848
R23431 VDD.n789 VDD.n675 749.848
R23432 VDD.n827 VDD.n675 749.848
R23433 VDD.n828 VDD.n827 749.848
R23434 VDD.n828 VDD.n669 749.848
R23435 VDD.n844 VDD.n669 749.848
R23436 VDD.n1183 VDD 516.447
R23437 VDD.n1191 VDD 475.642
R23438 VDD.n228 VDD.n227 293.12
R23439 VDD.n229 VDD.n228 293.12
R23440 VDD.n230 VDD.n229 293.12
R23441 VDD.n231 VDD.n230 293.12
R23442 VDD.n232 VDD.n231 293.12
R23443 VDD.t25 VDD.t31 264.177
R23444 VDD.t19 VDD.t25 264.177
R23445 VDD.t7 VDD.t19 264.177
R23446 VDD.t22 VDD.t28 264.177
R23447 VDD.t10 VDD.t22 264.177
R23448 VDD.t4 VDD.t1 264.177
R23449 VDD.t1 VDD.t16 264.177
R23450 VDD.t34 VDD.t13 264.177
R23451 VDD.n1526 VDD.n1525 259.666
R23452 VDD.n903 VDD.n902 259.666
R23453 VDD.n846 VDD.n845 259.666
R23454 VDD.n644 VDD.n643 259.666
R23455 VDD.n623 VDD.n622 259.666
R23456 VDD.n1186 VDD.n188 259.666
R23457 VDD.n1179 VDD.n191 259.666
R23458 VDD.n245 VDD.t33 222.22
R23459 VDD.n1520 VDD.n1519 185
R23460 VDD.n1512 VDD.n1511 185
R23461 VDD.n1501 VDD.n1500 185
R23462 VDD.n1493 VDD.n1492 185
R23463 VDD.n1485 VDD.n1484 185
R23464 VDD.n1306 VDD.n1305 185
R23465 VDD.n1316 VDD.n1315 185
R23466 VDD.n1324 VDD.n1323 185
R23467 VDD.n1332 VDD.n1331 185
R23468 VDD.n1340 VDD.n1339 185
R23469 VDD.n1350 VDD.n1349 185
R23470 VDD.n1358 VDD.n1357 185
R23471 VDD.n1366 VDD.n1365 185
R23472 VDD.n1374 VDD.n1373 185
R23473 VDD.n1384 VDD.n1383 185
R23474 VDD.n1392 VDD.n1391 185
R23475 VDD.n1400 VDD.n1399 185
R23476 VDD.n1408 VDD.n1407 185
R23477 VDD.n1418 VDD.n1417 185
R23478 VDD.n901 VDD.n900 185
R23479 VDD.n892 VDD.n870 185
R23480 VDD.n844 VDD.n843 185
R23481 VDD.n836 VDD.n669 185
R23482 VDD.n829 VDD.n828 185
R23483 VDD.n827 VDD.n826 185
R23484 VDD.n679 VDD.n675 185
R23485 VDD.n789 VDD.n681 185
R23486 VDD.n790 VDD.n683 185
R23487 VDD.n791 VDD.n685 185
R23488 VDD.n793 VDD.n792 185
R23489 VDD.n788 VDD.n787 185
R23490 VDD.n780 VDD.n690 185
R23491 VDD.n774 VDD.n773 185
R23492 VDD.n772 VDD.n771 185
R23493 VDD.n761 VDD.n696 185
R23494 VDD.n755 VDD.n754 185
R23495 VDD.n753 VDD.n752 185
R23496 VDD.n707 VDD.n703 185
R23497 VDD.n713 VDD.n709 185
R23498 VDD.n714 VDD.n711 185
R23499 VDD.n642 VDD.n641 185
R23500 VDD.n634 VDD.n633 185
R23501 VDD.n632 VDD.n631 185
R23502 VDD.n617 VDD.n616 185
R23503 VDD.n609 VDD.n608 185
R23504 VDD.n599 VDD.n598 185
R23505 VDD.n591 VDD.n590 185
R23506 VDD.n582 VDD.n581 185
R23507 VDD.n574 VDD.n573 185
R23508 VDD.n564 VDD.n563 185
R23509 VDD.n556 VDD.n555 185
R23510 VDD.n548 VDD.n547 185
R23511 VDD.n540 VDD.n539 185
R23512 VDD.n530 VDD.n529 185
R23513 VDD.n522 VDD.n521 185
R23514 VDD.n514 VDD.n513 185
R23515 VDD.n506 VDD.n505 185
R23516 VDD.n496 VDD.n495 185
R23517 VDD.n488 VDD.n487 185
R23518 VDD.n480 VDD.n479 185
R23519 VDD.n472 VDD.n471 185
R23520 VDD.n462 VDD.n461 185
R23521 VDD.t13 VDD.n642 178.233
R23522 VDD.n366 VDD.n365 176.62
R23523 VDD.n632 VDD.t7 171.311
R23524 VDD.n253 VDD.t3 166.1
R23525 VDD.n251 VDD.t0 166.1
R23526 VDD.n242 VDD.t9 166.1
R23527 VDD.n244 VDD.t15 166.1
R23528 VDD.n241 VDD.t21 166.1
R23529 VDD.n246 VDD.t12 166.1
R23530 VDD.n260 VDD.t27 166.1
R23531 VDD.n262 VDD.t6 166.099
R23532 VDD.n239 VDD.t18 166.098
R23533 VDD.n267 VDD.t24 166.098
R23534 VDD.n269 VDD.t30 166.097
R23535 VDD.n242 VDD.n241 161.952
R23536 VDD.n254 VDD.n242 154.24
R23537 VDD.n227 VDD 147.84
R23538 VDD.n259 VDD.n241 146.528
R23539 VDD.n633 VDD.t4 135.549
R23540 VDD.n633 VDD.t10 128.627
R23541 VDD.n253 VDD.n252 127.248
R23542 VDD.n269 VDD.n268 123.392
R23543 VDD.n248 VDD.n245 122.204
R23544 VDD.n261 VDD.n260 119.536
R23545 VDD.n646 VDD.n232 110.136
R23546 VDD.n251 VDD.n250 100.256
R23547 VDD.n267 VDD.n266 96.4
R23548 VDD.t28 VDD.n632 92.865
R23549 VDD.n263 VDD.n262 92.544
R23550 VDD.n1192 VDD.n185 89.734
R23551 VDD.n247 VDD.n246 88.688
R23552 VDD.n270 VDD.n269 87.568
R23553 VDD.n642 VDD.t16 85.944
R23554 VDD.n903 VDD.n869 85.333
R23555 VDD.n894 VDD.n893 85.333
R23556 VDD.n894 VDD.n871 85.333
R23557 VDD.n887 VDD.n873 85.333
R23558 VDD.n891 VDD.n873 85.333
R23559 VDD.n846 VDD.n668 85.333
R23560 VDD.n838 VDD.n837 85.333
R23561 VDD.n838 VDD.n670 85.333
R23562 VDD.n830 VDD.n672 85.333
R23563 VDD.n835 VDD.n672 85.333
R23564 VDD.n825 VDD.n677 85.333
R23565 VDD.n677 VDD.n674 85.333
R23566 VDD.n820 VDD.n819 85.333
R23567 VDD.n814 VDD.n813 85.333
R23568 VDD.n815 VDD.n814 85.333
R23569 VDD.n809 VDD.n808 85.333
R23570 VDD.n810 VDD.n809 85.333
R23571 VDD.n804 VDD.n803 85.333
R23572 VDD.n805 VDD.n804 85.333
R23573 VDD.n799 VDD.n798 85.333
R23574 VDD.n786 VDD.n689 85.333
R23575 VDD.n794 VDD.n689 85.333
R23576 VDD.n782 VDD.n781 85.333
R23577 VDD.n782 VDD.n691 85.333
R23578 VDD.n775 VDD.n693 85.333
R23579 VDD.n779 VDD.n693 85.333
R23580 VDD.n766 VDD.n698 85.333
R23581 VDD.n763 VDD.n762 85.333
R23582 VDD.n763 VDD.n697 85.333
R23583 VDD.n756 VDD.n700 85.333
R23584 VDD.n760 VDD.n700 85.333
R23585 VDD.n751 VDD.n705 85.333
R23586 VDD.n705 VDD.n702 85.333
R23587 VDD.n746 VDD.n745 85.333
R23588 VDD.n740 VDD.n739 85.333
R23589 VDD.n741 VDD.n740 85.333
R23590 VDD.n735 VDD.n734 85.333
R23591 VDD.n736 VDD.n735 85.333
R23592 VDD.n730 VDD.n729 85.333
R23593 VDD.n731 VDD.n730 85.333
R23594 VDD.n644 VDD.n234 85.333
R23595 VDD.n636 VDD.n635 85.333
R23596 VDD.n636 VDD.n235 85.333
R23597 VDD.n630 VDD.n626 85.333
R23598 VDD.n626 VDD.n237 85.333
R23599 VDD.n270 VDD.n238 85.333
R23600 VDD.n265 VDD.n238 85.333
R23601 VDD.n265 VDD.n264 85.333
R23602 VDD.n264 VDD.n240 85.333
R23603 VDD.n258 VDD.n240 85.333
R23604 VDD.n258 VDD.n257 85.333
R23605 VDD.n257 VDD.n256 85.333
R23606 VDD.n256 VDD.n255 85.333
R23607 VDD.n255 VDD.n243 85.333
R23608 VDD.n249 VDD.n243 85.333
R23609 VDD.n249 VDD.n248 85.333
R23610 VDD.n1187 VDD.n1186 85.333
R23611 VDD.n1180 VDD.n1179 85.333
R23612 VDD.n899 VDD.n869 82.651
R23613 VDD.n842 VDD.n668 82.651
R23614 VDD.n819 VDD.n818 82.651
R23615 VDD.n798 VDD.n687 82.651
R23616 VDD.n770 VDD.n698 82.651
R23617 VDD.n745 VDD.n744 82.651
R23618 VDD.n640 VDD.n234 82.651
R23619 VDD.n1188 VDD.n1187 82.651
R23620 VDD.n1181 VDD.n1180 82.651
R23621 VDD.n820 VDD.n676 80.7
R23622 VDD.n800 VDD.n799 80.7
R23623 VDD.n766 VDD.n695 80.7
R23624 VDD.n746 VDD.n704 80.7
R23625 VDD.n268 VDD.n238 76
R23626 VDD.n257 VDD.n241 76
R23627 VDD.n256 VDD.n242 76
R23628 VDD.n266 VDD.n265 76
R23629 VDD.n264 VDD.n263 76
R23630 VDD.n261 VDD.n240 76
R23631 VDD.n259 VDD.n258 76
R23632 VDD.n255 VDD.n254 76
R23633 VDD.n252 VDD.n243 76
R23634 VDD.n250 VDD.n249 76
R23635 VDD.n248 VDD.n247 76
R23636 VDD.n247 VDD.n244 73.264
R23637 VDD.n246 VDD.n245 69.888
R23638 VDD.n263 VDD.n239 69.408
R23639 VDD.n1184 VDD.n189 67.425
R23640 VDD.n826 VDD.n825 66.803
R23641 VDD.n803 VDD.n685 66.803
R23642 VDD.n775 VDD.n774 66.803
R23643 VDD.n752 VDD.n751 66.803
R23644 VDD.n729 VDD.n715 66.803
R23645 VDD.n266 VDD.n239 65.552
R23646 VDD.n900 VDD.n871 63.024
R23647 VDD.n843 VDD.n670 63.024
R23648 VDD.n815 VDD.n679 63.024
R23649 VDD.n794 VDD.n793 63.024
R23650 VDD.n771 VDD.n697 63.024
R23651 VDD.n741 VDD.n707 63.024
R23652 VDD.n641 VDD.n235 63.024
R23653 VDD.n187 VDD.n185 63.024
R23654 VDD.n250 VDD.n244 61.696
R23655 VDD.n366 VDD.n364 54.344
R23656 VDD.n349 VDD.n348 54.344
R23657 VDD.n377 VDD.n376 47.551
R23658 VDD.n338 VDD.n337 47.551
R23659 VDD.n887 VDD.n886 45.47
R23660 VDD.n830 VDD.n829 45.47
R23661 VDD.n808 VDD.n683 45.47
R23662 VDD.n781 VDD.n780 45.47
R23663 VDD.n756 VDD.n755 45.47
R23664 VDD.n734 VDD.n711 45.47
R23665 VDD.n631 VDD.n630 45.47
R23666 VDD.n431 VDD.n430 44.155
R23667 VDD.n282 VDD.n281 44.155
R23668 VDD.n262 VDD.n261 42.416
R23669 VDD.n892 VDD.n891 41.691
R23670 VDD.n836 VDD.n835 41.691
R23671 VDD.n810 VDD.n681 41.691
R23672 VDD.n787 VDD.n691 41.691
R23673 VDD.n761 VDD.n760 41.691
R23674 VDD.n736 VDD.n709 41.691
R23675 VDD.n634 VDD.n237 41.691
R23676 VDD.n388 VDD.n387 40.758
R23677 VDD.n327 VDD.n326 40.758
R23678 VDD.n268 VDD.n267 38.56
R23679 VDD.n420 VDD.n419 37.362
R23680 VDD.n293 VDD.n292 37.362
R23681 VDD VDD.n270 34.986
R23682 VDD.n252 VDD.n251 34.704
R23683 VDD.n589 VDD.n443 34.216
R23684 VDD.n399 VDD.n398 33.965
R23685 VDD.n316 VDD.n315 33.965
R23686 VDD.n232 VDD.n221 32.824
R23687 VDD.n231 VDD.n222 32.824
R23688 VDD.n230 VDD.n223 32.824
R23689 VDD.n229 VDD.n224 32.824
R23690 VDD.n228 VDD.n225 32.824
R23691 VDD.n227 VDD.n226 32.824
R23692 VDD.n409 VDD.n408 30.568
R23693 VDD.n304 VDD.n303 30.568
R23694 VDD.n410 VDD.n409 27.172
R23695 VDD.n305 VDD.n304 27.172
R23696 VDD.n271 VDD 26.186
R23697 VDD.n1068 VDD 24.8
R23698 VDD.n886 VDD.n885 24.758
R23699 VDD.n631 VDD.n625 24.758
R23700 VDD.n1513 VDD.n1512 24.137
R23701 VDD.n1307 VDD.n1306 24.137
R23702 VDD.n1341 VDD.n1340 24.137
R23703 VDD.n1375 VDD.n1374 24.137
R23704 VDD.n1409 VDD.n1408 24.137
R23705 VDD.n893 VDD.n892 24.137
R23706 VDD.n837 VDD.n836 24.137
R23707 VDD.n813 VDD.n681 24.137
R23708 VDD.n787 VDD.n786 24.137
R23709 VDD.n762 VDD.n761 24.137
R23710 VDD.n739 VDD.n709 24.137
R23711 VDD.n635 VDD.n634 24.137
R23712 VDD.n610 VDD.n609 24.137
R23713 VDD.n575 VDD.n574 24.137
R23714 VDD.n541 VDD.n540 24.137
R23715 VDD.n507 VDD.n506 24.137
R23716 VDD.n473 VDD.n472 24.137
R23717 VDD.n398 VDD.n397 23.775
R23718 VDD.n315 VDD.n314 23.775
R23719 VDD.n1037 VDD 21.329
R23720 VDD.n1450 VDD 21.072
R23721 VDD.n421 VDD.n420 20.379
R23722 VDD.n294 VDD.n293 20.379
R23723 VDD.n1502 VDD.n1501 20.357
R23724 VDD.n1317 VDD.n1316 20.357
R23725 VDD.n1351 VDD.n1350 20.357
R23726 VDD.n1385 VDD.n1384 20.357
R23727 VDD.n1419 VDD.n1418 20.357
R23728 VDD.n829 VDD.n674 20.357
R23729 VDD.n805 VDD.n683 20.357
R23730 VDD.n780 VDD.n779 20.357
R23731 VDD.n755 VDD.n702 20.357
R23732 VDD.n731 VDD.n711 20.357
R23733 VDD.n600 VDD.n599 20.357
R23734 VDD.n565 VDD.n564 20.357
R23735 VDD.n531 VDD.n530 20.357
R23736 VDD.n497 VDD.n496 20.357
R23737 VDD.n463 VDD.n462 20.357
R23738 VDD.n1005 VDD 18.47
R23739 VDD.n1529 VDD.n1527 17.81
R23740 VDD.n387 VDD.n386 16.982
R23741 VDD.n326 VDD.n325 16.982
R23742 VDD.n974 VDD 15.612
R23743 VDD.n260 VDD.n259 15.424
R23744 VDD.n432 VDD.n431 13.586
R23745 VDD.n283 VDD.n282 13.586
R23746 VDD VDD.n1004 13.313
R23747 VDD VDD.n973 13.313
R23748 VDD VDD.n884 13.313
R23749 VDD VDD.n936 13.313
R23750 VDD.n357 VDD.n356 13.176
R23751 VDD.n942 VDD 10.814
R23752 VDD.n376 VDD.n375 10.189
R23753 VDD.n337 VDD.n336 10.189
R23754 VDD.n438 VDD.n437 9.3
R23755 VDD.n427 VDD.n426 9.3
R23756 VDD.n416 VDD.n415 9.3
R23757 VDD.n405 VDD.n404 9.3
R23758 VDD.n394 VDD.n393 9.3
R23759 VDD.n383 VDD.n382 9.3
R23760 VDD.n372 VDD.n371 9.3
R23761 VDD.n360 VDD.n359 9.3
R23762 VDD.n353 VDD.n352 9.3
R23763 VDD.n342 VDD.n341 9.3
R23764 VDD.n331 VDD.n330 9.3
R23765 VDD.n320 VDD.n319 9.3
R23766 VDD.n309 VDD.n308 9.3
R23767 VDD.n298 VDD.n297 9.3
R23768 VDD.n287 VDD.n286 9.3
R23769 VDD.n276 VDD.n275 9.3
R23770 VDD.n274 VDD.n273 9.3
R23771 VDD.n278 VDD.n277 9.3
R23772 VDD.n285 VDD.n284 9.3
R23773 VDD.n284 VDD.n283 9.3
R23774 VDD.n289 VDD.n288 9.3
R23775 VDD.n296 VDD.n295 9.3
R23776 VDD.n295 VDD.n294 9.3
R23777 VDD.n300 VDD.n299 9.3
R23778 VDD.n307 VDD.n306 9.3
R23779 VDD.n306 VDD.n305 9.3
R23780 VDD.n311 VDD.n310 9.3
R23781 VDD.n318 VDD.n317 9.3
R23782 VDD.n317 VDD.n316 9.3
R23783 VDD.n322 VDD.n321 9.3
R23784 VDD.n329 VDD.n328 9.3
R23785 VDD.n328 VDD.n327 9.3
R23786 VDD.n333 VDD.n332 9.3
R23787 VDD.n340 VDD.n339 9.3
R23788 VDD.n339 VDD.n338 9.3
R23789 VDD.n344 VDD.n343 9.3
R23790 VDD.n351 VDD.n350 9.3
R23791 VDD.n350 VDD.n349 9.3
R23792 VDD.n355 VDD.n354 9.3
R23793 VDD.n358 VDD.n357 9.3
R23794 VDD.n368 VDD.n367 9.3
R23795 VDD.n367 VDD.n366 9.3
R23796 VDD.n370 VDD.n369 9.3
R23797 VDD.n379 VDD.n378 9.3
R23798 VDD.n378 VDD.n377 9.3
R23799 VDD.n381 VDD.n380 9.3
R23800 VDD.n390 VDD.n389 9.3
R23801 VDD.n389 VDD.n388 9.3
R23802 VDD.n392 VDD.n391 9.3
R23803 VDD.n401 VDD.n400 9.3
R23804 VDD.n400 VDD.n399 9.3
R23805 VDD.n403 VDD.n402 9.3
R23806 VDD.n412 VDD.n411 9.3
R23807 VDD.n411 VDD.n410 9.3
R23808 VDD.n414 VDD.n413 9.3
R23809 VDD.n423 VDD.n422 9.3
R23810 VDD.n422 VDD.n421 9.3
R23811 VDD.n425 VDD.n424 9.3
R23812 VDD.n434 VDD.n433 9.3
R23813 VDD.n433 VDD.n432 9.3
R23814 VDD.n436 VDD.n435 9.3
R23815 VDD.n441 VDD.n440 9.3
R23816 VDD VDD.n847 8.141
R23817 VDD.n1425 VDD.n1302 8.045
R23818 VDD.n727 VDD.n715 8.045
R23819 VDD.n456 VDD.n455 8.045
R23820 VDD VDD.n646 8.032
R23821 VDD.n254 VDD.n253 7.712
R23822 VDD VDD.n1067 6.334
R23823 VDD VDD.n1448 6.26
R23824 VDD.n367 VDD.n362 6.023
R23825 VDD.n350 VDD.n346 6.023
R23826 VDD.n940 VDD 5.855
R23827 VDD VDD.n941 5.744
R23828 VDD.n941 VDD 5.542
R23829 VDD.n1521 VDD.n1520 5.485
R23830 VDD.n1486 VDD.n1485 5.485
R23831 VDD.n1333 VDD.n1332 5.485
R23832 VDD.n1367 VDD.n1366 5.485
R23833 VDD.n1401 VDD.n1400 5.485
R23834 VDD.n900 VDD.n899 5.485
R23835 VDD.n843 VDD.n842 5.485
R23836 VDD.n818 VDD.n679 5.485
R23837 VDD.n793 VDD.n687 5.485
R23838 VDD.n771 VDD.n770 5.485
R23839 VDD.n744 VDD.n707 5.485
R23840 VDD.n641 VDD.n640 5.485
R23841 VDD.n618 VDD.n617 5.485
R23842 VDD.n583 VDD.n582 5.485
R23843 VDD.n549 VDD.n548 5.485
R23844 VDD.n515 VDD.n514 5.485
R23845 VDD.n481 VDD.n480 5.485
R23846 VDD.n1188 VDD.n187 5.485
R23847 VDD.n1181 VDD.n189 5.485
R23848 VDD.n378 VDD.n374 5.27
R23849 VDD.n339 VDD.n335 5.27
R23850 VDD.n429 VDD.n428 4.894
R23851 VDD.n280 VDD.n279 4.894
R23852 VDD.n442 VDD.n441 4.84
R23853 VDD.n888 VDD.n887 4.65
R23854 VDD.n889 VDD.n873 4.65
R23855 VDD.n891 VDD.n890 4.65
R23856 VDD.n893 VDD.n872 4.65
R23857 VDD.n895 VDD.n894 4.65
R23858 VDD.n896 VDD.n871 4.65
R23859 VDD.n899 VDD.n898 4.65
R23860 VDD.n897 VDD.n869 4.65
R23861 VDD.n904 VDD.n903 4.65
R23862 VDD.n729 VDD.n728 4.65
R23863 VDD.n730 VDD.n712 4.65
R23864 VDD.n732 VDD.n731 4.65
R23865 VDD.n734 VDD.n733 4.65
R23866 VDD.n735 VDD.n710 4.65
R23867 VDD.n737 VDD.n736 4.65
R23868 VDD.n739 VDD.n738 4.65
R23869 VDD.n740 VDD.n708 4.65
R23870 VDD.n742 VDD.n741 4.65
R23871 VDD.n744 VDD.n743 4.65
R23872 VDD.n745 VDD.n706 4.65
R23873 VDD.n747 VDD.n746 4.65
R23874 VDD.n748 VDD.n704 4.65
R23875 VDD.n751 VDD.n750 4.65
R23876 VDD.n749 VDD.n705 4.65
R23877 VDD.n702 VDD.n701 4.65
R23878 VDD.n757 VDD.n756 4.65
R23879 VDD.n758 VDD.n700 4.65
R23880 VDD.n760 VDD.n759 4.65
R23881 VDD.n762 VDD.n699 4.65
R23882 VDD.n764 VDD.n763 4.65
R23883 VDD.n765 VDD.n697 4.65
R23884 VDD.n770 VDD.n769 4.65
R23885 VDD.n768 VDD.n698 4.65
R23886 VDD.n767 VDD.n766 4.65
R23887 VDD.n695 VDD.n694 4.65
R23888 VDD.n776 VDD.n775 4.65
R23889 VDD.n777 VDD.n693 4.65
R23890 VDD.n779 VDD.n778 4.65
R23891 VDD.n781 VDD.n692 4.65
R23892 VDD.n783 VDD.n782 4.65
R23893 VDD.n784 VDD.n691 4.65
R23894 VDD.n786 VDD.n785 4.65
R23895 VDD.n689 VDD.n688 4.65
R23896 VDD.n795 VDD.n794 4.65
R23897 VDD.n796 VDD.n687 4.65
R23898 VDD.n798 VDD.n797 4.65
R23899 VDD.n799 VDD.n686 4.65
R23900 VDD.n801 VDD.n800 4.65
R23901 VDD.n803 VDD.n802 4.65
R23902 VDD.n804 VDD.n684 4.65
R23903 VDD.n806 VDD.n805 4.65
R23904 VDD.n808 VDD.n807 4.65
R23905 VDD.n809 VDD.n682 4.65
R23906 VDD.n811 VDD.n810 4.65
R23907 VDD.n813 VDD.n812 4.65
R23908 VDD.n814 VDD.n680 4.65
R23909 VDD.n816 VDD.n815 4.65
R23910 VDD.n818 VDD.n817 4.65
R23911 VDD.n819 VDD.n678 4.65
R23912 VDD.n821 VDD.n820 4.65
R23913 VDD.n822 VDD.n676 4.65
R23914 VDD.n825 VDD.n824 4.65
R23915 VDD.n823 VDD.n677 4.65
R23916 VDD.n674 VDD.n673 4.65
R23917 VDD.n831 VDD.n830 4.65
R23918 VDD.n833 VDD.n672 4.65
R23919 VDD.n835 VDD.n834 4.65
R23920 VDD.n837 VDD.n671 4.65
R23921 VDD.n839 VDD.n838 4.65
R23922 VDD.n840 VDD.n670 4.65
R23923 VDD.n842 VDD.n841 4.65
R23924 VDD.n668 VDD.n667 4.65
R23925 VDD.n847 VDD.n846 4.65
R23926 VDD.n458 VDD.n457 4.65
R23927 VDD.n460 VDD.n459 4.65
R23928 VDD.n464 VDD.n463 4.65
R23929 VDD.n466 VDD.n465 4.65
R23930 VDD.n468 VDD.n467 4.65
R23931 VDD.n470 VDD.n469 4.65
R23932 VDD.n474 VDD.n473 4.65
R23933 VDD.n476 VDD.n475 4.65
R23934 VDD.n478 VDD.n477 4.65
R23935 VDD.n482 VDD.n481 4.65
R23936 VDD.n484 VDD.n483 4.65
R23937 VDD.n486 VDD.n485 4.65
R23938 VDD.n490 VDD.n489 4.65
R23939 VDD.n492 VDD.n491 4.65
R23940 VDD.n494 VDD.n493 4.65
R23941 VDD.n498 VDD.n497 4.65
R23942 VDD.n500 VDD.n499 4.65
R23943 VDD.n502 VDD.n501 4.65
R23944 VDD.n504 VDD.n503 4.65
R23945 VDD.n508 VDD.n507 4.65
R23946 VDD.n510 VDD.n509 4.65
R23947 VDD.n512 VDD.n511 4.65
R23948 VDD.n516 VDD.n515 4.65
R23949 VDD.n518 VDD.n517 4.65
R23950 VDD.n520 VDD.n519 4.65
R23951 VDD.n524 VDD.n523 4.65
R23952 VDD.n526 VDD.n525 4.65
R23953 VDD.n528 VDD.n527 4.65
R23954 VDD.n532 VDD.n531 4.65
R23955 VDD.n534 VDD.n533 4.65
R23956 VDD.n536 VDD.n535 4.65
R23957 VDD.n538 VDD.n537 4.65
R23958 VDD.n542 VDD.n541 4.65
R23959 VDD.n544 VDD.n543 4.65
R23960 VDD.n546 VDD.n545 4.65
R23961 VDD.n550 VDD.n549 4.65
R23962 VDD.n552 VDD.n551 4.65
R23963 VDD.n554 VDD.n553 4.65
R23964 VDD.n558 VDD.n557 4.65
R23965 VDD.n560 VDD.n559 4.65
R23966 VDD.n562 VDD.n561 4.65
R23967 VDD.n566 VDD.n565 4.65
R23968 VDD.n568 VDD.n567 4.65
R23969 VDD.n570 VDD.n569 4.65
R23970 VDD.n572 VDD.n571 4.65
R23971 VDD.n576 VDD.n575 4.65
R23972 VDD.n578 VDD.n577 4.65
R23973 VDD.n580 VDD.n579 4.65
R23974 VDD.n584 VDD.n583 4.65
R23975 VDD.n586 VDD.n585 4.65
R23976 VDD.n588 VDD.n587 4.65
R23977 VDD.n593 VDD.n592 4.65
R23978 VDD.n595 VDD.n594 4.65
R23979 VDD.n597 VDD.n596 4.65
R23980 VDD.n601 VDD.n600 4.65
R23981 VDD.n603 VDD.n602 4.65
R23982 VDD.n605 VDD.n604 4.65
R23983 VDD.n607 VDD.n606 4.65
R23984 VDD.n611 VDD.n610 4.65
R23985 VDD.n613 VDD.n612 4.65
R23986 VDD.n615 VDD.n614 4.65
R23987 VDD.n619 VDD.n618 4.65
R23988 VDD.n621 VDD.n620 4.65
R23989 VDD.n624 VDD.n623 4.65
R23990 VDD.n630 VDD.n629 4.65
R23991 VDD.n628 VDD.n626 4.65
R23992 VDD.n627 VDD.n237 4.65
R23993 VDD.n635 VDD.n236 4.65
R23994 VDD.n637 VDD.n636 4.65
R23995 VDD.n638 VDD.n235 4.65
R23996 VDD.n640 VDD.n639 4.65
R23997 VDD.n234 VDD.n233 4.65
R23998 VDD.n645 VDD.n644 4.65
R23999 VDD.n1190 VDD.n185 4.65
R24000 VDD.n1189 VDD.n1188 4.65
R24001 VDD.n1187 VDD.n186 4.65
R24002 VDD.n1186 VDD.n1185 4.65
R24003 VDD.n1182 VDD.n1181 4.65
R24004 VDD.n1180 VDD.n190 4.65
R24005 VDD.n1179 VDD.n1178 4.65
R24006 VDD.n1424 VDD.n1423 4.65
R24007 VDD.n1422 VDD.n1421 4.65
R24008 VDD.n1420 VDD.n1419 4.65
R24009 VDD.n1416 VDD.n1415 4.65
R24010 VDD.n1414 VDD.n1413 4.65
R24011 VDD.n1412 VDD.n1411 4.65
R24012 VDD.n1410 VDD.n1409 4.65
R24013 VDD.n1406 VDD.n1405 4.65
R24014 VDD.n1404 VDD.n1403 4.65
R24015 VDD.n1402 VDD.n1401 4.65
R24016 VDD.n1398 VDD.n1397 4.65
R24017 VDD.n1396 VDD.n1395 4.65
R24018 VDD.n1394 VDD.n1393 4.65
R24019 VDD.n1390 VDD.n1389 4.65
R24020 VDD.n1388 VDD.n1387 4.65
R24021 VDD.n1386 VDD.n1385 4.65
R24022 VDD.n1382 VDD.n1381 4.65
R24023 VDD.n1380 VDD.n1379 4.65
R24024 VDD.n1378 VDD.n1377 4.65
R24025 VDD.n1376 VDD.n1375 4.65
R24026 VDD.n1372 VDD.n1371 4.65
R24027 VDD.n1370 VDD.n1369 4.65
R24028 VDD.n1368 VDD.n1367 4.65
R24029 VDD.n1364 VDD.n1363 4.65
R24030 VDD.n1362 VDD.n1361 4.65
R24031 VDD.n1360 VDD.n1359 4.65
R24032 VDD.n1356 VDD.n1355 4.65
R24033 VDD.n1354 VDD.n1353 4.65
R24034 VDD.n1352 VDD.n1351 4.65
R24035 VDD.n1348 VDD.n1347 4.65
R24036 VDD.n1346 VDD.n1345 4.65
R24037 VDD.n1344 VDD.n1343 4.65
R24038 VDD.n1342 VDD.n1341 4.65
R24039 VDD.n1338 VDD.n1337 4.65
R24040 VDD.n1336 VDD.n1335 4.65
R24041 VDD.n1334 VDD.n1333 4.65
R24042 VDD.n1330 VDD.n1329 4.65
R24043 VDD.n1328 VDD.n1327 4.65
R24044 VDD.n1326 VDD.n1325 4.65
R24045 VDD.n1322 VDD.n1321 4.65
R24046 VDD.n1320 VDD.n1319 4.65
R24047 VDD.n1318 VDD.n1317 4.65
R24048 VDD.n1314 VDD.n1313 4.65
R24049 VDD.n1312 VDD.n1311 4.65
R24050 VDD.n1310 VDD.n1309 4.65
R24051 VDD.n1308 VDD.n1307 4.65
R24052 VDD.n1304 VDD.n1303 4.65
R24053 VDD.n1483 VDD.n1482 4.65
R24054 VDD.n1487 VDD.n1486 4.65
R24055 VDD.n1489 VDD.n1488 4.65
R24056 VDD.n1491 VDD.n1490 4.65
R24057 VDD.n1495 VDD.n1494 4.65
R24058 VDD.n1497 VDD.n1496 4.65
R24059 VDD.n1499 VDD.n1498 4.65
R24060 VDD.n1503 VDD.n1502 4.65
R24061 VDD.n1505 VDD.n1504 4.65
R24062 VDD.n1508 VDD.n1507 4.65
R24063 VDD.n1510 VDD.n1509 4.65
R24064 VDD.n1514 VDD.n1513 4.65
R24065 VDD.n1516 VDD.n1515 4.65
R24066 VDD.n1518 VDD.n1517 4.65
R24067 VDD.n1522 VDD.n1521 4.65
R24068 VDD.n1524 VDD.n1523 4.65
R24069 VDD.n1527 VDD.n1526 4.65
R24070 VDD.n389 VDD.n385 4.517
R24071 VDD.n328 VDD.n324 4.517
R24072 VDD VDD.n1036 4.497
R24073 VDD VDD.n726 4.497
R24074 VDD.n1193 VDD 4.497
R24075 VDD.n221 VDD.t14 4.428
R24076 VDD.n221 VDD.t35 4.428
R24077 VDD.n222 VDD.t2 4.428
R24078 VDD.n222 VDD.t17 4.428
R24079 VDD.n223 VDD.t11 4.428
R24080 VDD.n223 VDD.t5 4.428
R24081 VDD.n224 VDD.t29 4.428
R24082 VDD.n224 VDD.t23 4.428
R24083 VDD.n225 VDD.t20 4.428
R24084 VDD.n225 VDD.t8 4.428
R24085 VDD.n226 VDD.t32 4.428
R24086 VDD.n226 VDD.t26 4.428
R24087 VDD.n940 VDD.n939 4.372
R24088 VDD VDD.n904 4.339
R24089 VDD.n937 VDD 4.273
R24090 VDD.n418 VDD.n417 4.141
R24091 VDD.n291 VDD.n290 4.141
R24092 VDD.n456 VDD.n454 3.781
R24093 VDD.n400 VDD.n396 3.764
R24094 VDD.n317 VDD.n313 3.764
R24095 VDD.n1185 VDD 3.723
R24096 VDD.n1426 VDD.n1425 3.707
R24097 VDD.n1494 VDD.n1493 3.657
R24098 VDD.n1325 VDD.n1324 3.657
R24099 VDD.n1359 VDD.n1358 3.657
R24100 VDD.n1393 VDD.n1392 3.657
R24101 VDD.n826 VDD.n676 3.657
R24102 VDD.n800 VDD.n685 3.657
R24103 VDD.n774 VDD.n695 3.657
R24104 VDD.n752 VDD.n704 3.657
R24105 VDD.n592 VDD.n591 3.657
R24106 VDD.n557 VDD.n556 3.657
R24107 VDD.n523 VDD.n522 3.657
R24108 VDD.n489 VDD.n488 3.657
R24109 VDD.n364 VDD.n363 3.396
R24110 VDD.n348 VDD.n347 3.396
R24111 VDD.n407 VDD.n406 3.388
R24112 VDD.n302 VDD.n301 3.388
R24113 VDD.n727 VDD 3.16
R24114 VDD.n939 VDD.n938 3.089
R24115 VDD.n411 VDD.n407 3.011
R24116 VDD.n306 VDD.n302 3.011
R24117 VDD.n938 VDD.n937 2.913
R24118 VDD.n905 VDD 2.904
R24119 VDD.n848 VDD 2.904
R24120 VDD VDD.n1177 2.904
R24121 VDD.n396 VDD.n395 2.635
R24122 VDD.n313 VDD.n312 2.635
R24123 VDD.n647 VDD 2.495
R24124 VDD.n625 VDD 2.343
R24125 VDD.n422 VDD.n418 2.258
R24126 VDD.n295 VDD.n291 2.258
R24127 VDD.n885 VDD 2.139
R24128 VDD VDD.n940 2.026
R24129 VDD.n941 VDD 1.985
R24130 VDD VDD.n1184 1.884
R24131 VDD.n385 VDD.n384 1.882
R24132 VDD.n324 VDD.n323 1.882
R24133 VDD.n1561 VDD.n0 1.7
R24134 VDD.n194 VDD.n193 1.7
R24135 VDD.n433 VDD.n429 1.505
R24136 VDD.n284 VDD.n280 1.505
R24137 VDD VDD.n1192 1.419
R24138 VDD.n937 VDD 1.22
R24139 VDD.n938 VDD 1.22
R24140 VDD.n374 VDD.n373 1.129
R24141 VDD.n335 VDD.n334 1.129
R24142 VDD VDD.n624 1.126
R24143 VDD.n1178 VDD 1.126
R24144 VDD.n939 VDD 1.045
R24145 VDD.n1084 VDD.n1083 0.852
R24146 VDD.n1084 VDD.n1078 0.852
R24147 VDD.n1084 VDD.n1050 0.852
R24148 VDD.n1084 VDD.n1052 0.852
R24149 VDD.n1084 VDD.n1054 0.852
R24150 VDD.n1084 VDD.n1074 0.852
R24151 VDD.n1094 VDD.n1093 0.852
R24152 VDD.n1094 VDD.n1089 0.852
R24153 VDD.n1094 VDD.n1018 0.852
R24154 VDD.n1094 VDD.n1020 0.852
R24155 VDD.n1094 VDD.n1023 0.852
R24156 VDD.n1094 VDD.n1043 0.852
R24157 VDD.n1105 VDD.n1104 0.852
R24158 VDD.n1105 VDD.n1099 0.852
R24159 VDD.n1105 VDD.n987 0.852
R24160 VDD.n1105 VDD.n989 0.852
R24161 VDD.n1105 VDD.n991 0.852
R24162 VDD.n1105 VDD.n1011 0.852
R24163 VDD.n1115 VDD.n1114 0.852
R24164 VDD.n1115 VDD.n1110 0.852
R24165 VDD.n1115 VDD.n955 0.852
R24166 VDD.n1115 VDD.n957 0.852
R24167 VDD.n1115 VDD.n960 0.852
R24168 VDD.n1115 VDD.n980 0.852
R24169 VDD.n1125 VDD.n1124 0.852
R24170 VDD.n1125 VDD.n1120 0.852
R24171 VDD.n1125 VDD.n918 0.852
R24172 VDD.n1125 VDD.n920 0.852
R24173 VDD.n1125 VDD.n923 0.852
R24174 VDD.n1125 VDD.n948 0.852
R24175 VDD.n1136 VDD.n1135 0.852
R24176 VDD.n1136 VDD.n1130 0.852
R24177 VDD.n1136 VDD.n861 0.852
R24178 VDD.n1136 VDD.n863 0.852
R24179 VDD.n1136 VDD.n865 0.852
R24180 VDD.n1136 VDD.n911 0.852
R24181 VDD.n1147 VDD.n1146 0.852
R24182 VDD.n1147 VDD.n1141 0.852
R24183 VDD.n1147 VDD.n660 0.852
R24184 VDD.n1147 VDD.n662 0.852
R24185 VDD.n1147 VDD.n664 0.852
R24186 VDD.n1147 VDD.n854 0.852
R24187 VDD.n1158 VDD.n1157 0.852
R24188 VDD.n1158 VDD.n1152 0.852
R24189 VDD.n1158 VDD.n214 0.852
R24190 VDD.n1158 VDD.n216 0.852
R24191 VDD.n1158 VDD.n218 0.852
R24192 VDD.n1158 VDD.n653 0.852
R24193 VDD.n1169 VDD.n1168 0.852
R24194 VDD.n1169 VDD.n1163 0.852
R24195 VDD.n1169 VDD.n203 0.852
R24196 VDD.n1169 VDD.n205 0.852
R24197 VDD.n1169 VDD.n207 0.852
R24198 VDD.n1170 VDD.n1169 0.852
R24199 VDD.n273 VDD.n272 0.851
R24200 VDD.n440 VDD.n439 0.851
R24201 VDD.n1084 VDD.n1081 0.849
R24202 VDD.n1094 VDD.n1091 0.849
R24203 VDD.n1105 VDD.n1102 0.849
R24204 VDD.n1115 VDD.n1112 0.849
R24205 VDD.n1125 VDD.n1122 0.849
R24206 VDD.n1136 VDD.n1133 0.849
R24207 VDD.n1147 VDD.n1144 0.849
R24208 VDD.n1158 VDD.n1155 0.849
R24209 VDD.n1169 VDD.n1166 0.849
R24210 VDD.n1558 VDD.n1557 0.849
R24211 VDD.n1558 VDD.n1549 0.849
R24212 VDD.n1558 VDD.n1547 0.849
R24213 VDD.n1558 VDD.n1544 0.849
R24214 VDD.n1558 VDD.n1542 0.849
R24215 VDD.n1558 VDD.n1539 0.849
R24216 VDD.n1558 VDD.n1537 0.849
R24217 VDD.n1437 VDD.n1273 0.849
R24218 VDD.n1437 VDD.n1264 0.849
R24219 VDD.n1437 VDD.n1262 0.849
R24220 VDD.n1437 VDD.n1259 0.849
R24221 VDD.n1437 VDD.n1257 0.849
R24222 VDD.n1437 VDD.n1254 0.849
R24223 VDD.n1438 VDD.n1437 0.849
R24224 VDD.n1208 VDD.n1207 0.677
R24225 VDD.n1477 VDD.n1476 0.677
R24226 VDD.n1213 VDD.n169 0.563
R24227 VDD.n1213 VDD.n167 0.563
R24228 VDD.n1213 VDD.n161 0.563
R24229 VDD.n1218 VDD.n148 0.563
R24230 VDD.n1218 VDD.n146 0.563
R24231 VDD.n1218 VDD.n140 0.563
R24232 VDD.n1223 VDD.n127 0.563
R24233 VDD.n1223 VDD.n125 0.563
R24234 VDD.n1223 VDD.n119 0.563
R24235 VDD.n1228 VDD.n106 0.563
R24236 VDD.n1228 VDD.n104 0.563
R24237 VDD.n1228 VDD.n98 0.563
R24238 VDD.n1233 VDD.n85 0.563
R24239 VDD.n1233 VDD.n83 0.563
R24240 VDD.n1233 VDD.n77 0.563
R24241 VDD.n1238 VDD.n64 0.563
R24242 VDD.n1238 VDD.n62 0.563
R24243 VDD.n1238 VDD.n56 0.563
R24244 VDD.n1243 VDD.n43 0.563
R24245 VDD.n1243 VDD.n41 0.563
R24246 VDD.n1243 VDD.n35 0.563
R24247 VDD.n1248 VDD.n22 0.563
R24248 VDD.n1248 VDD.n20 0.563
R24249 VDD.n1248 VDD.n14 0.563
R24250 VDD.n1432 VDD.n1285 0.563
R24251 VDD.n1432 VDD.n1290 0.563
R24252 VDD.n1432 VDD.n1295 0.563
R24253 VDD.n1432 VDD.n1431 0.563
R24254 VDD.n728 VDD.n727 0.439
R24255 VDD.n458 VDD.n456 0.439
R24256 VDD.n1425 VDD.n1424 0.439
R24257 VDD.n888 VDD.n885 0.438
R24258 VDD.n629 VDD.n625 0.438
R24259 VDD.n889 VDD.n888 0.416
R24260 VDD.n890 VDD.n889 0.416
R24261 VDD.n890 VDD.n872 0.416
R24262 VDD.n895 VDD.n872 0.416
R24263 VDD.n896 VDD.n895 0.416
R24264 VDD.n898 VDD.n896 0.416
R24265 VDD.n898 VDD.n897 0.416
R24266 VDD.n728 VDD.n712 0.416
R24267 VDD.n732 VDD.n712 0.416
R24268 VDD.n733 VDD.n732 0.416
R24269 VDD.n733 VDD.n710 0.416
R24270 VDD.n737 VDD.n710 0.416
R24271 VDD.n738 VDD.n737 0.416
R24272 VDD.n738 VDD.n708 0.416
R24273 VDD.n742 VDD.n708 0.416
R24274 VDD.n743 VDD.n742 0.416
R24275 VDD.n743 VDD.n706 0.416
R24276 VDD.n747 VDD.n706 0.416
R24277 VDD.n748 VDD.n747 0.416
R24278 VDD.n750 VDD.n748 0.416
R24279 VDD.n750 VDD.n749 0.416
R24280 VDD.n749 VDD.n701 0.416
R24281 VDD.n757 VDD.n701 0.416
R24282 VDD.n758 VDD.n757 0.416
R24283 VDD.n759 VDD.n758 0.416
R24284 VDD.n759 VDD.n699 0.416
R24285 VDD.n764 VDD.n699 0.416
R24286 VDD.n765 VDD.n764 0.416
R24287 VDD.n769 VDD.n765 0.416
R24288 VDD.n769 VDD.n768 0.416
R24289 VDD.n768 VDD.n767 0.416
R24290 VDD.n767 VDD.n694 0.416
R24291 VDD.n776 VDD.n694 0.416
R24292 VDD.n777 VDD.n776 0.416
R24293 VDD.n778 VDD.n777 0.416
R24294 VDD.n778 VDD.n692 0.416
R24295 VDD.n783 VDD.n692 0.416
R24296 VDD.n784 VDD.n783 0.416
R24297 VDD.n785 VDD.n784 0.416
R24298 VDD.n785 VDD.n688 0.416
R24299 VDD.n795 VDD.n688 0.416
R24300 VDD.n796 VDD.n795 0.416
R24301 VDD.n797 VDD.n796 0.416
R24302 VDD.n797 VDD.n686 0.416
R24303 VDD.n801 VDD.n686 0.416
R24304 VDD.n802 VDD.n801 0.416
R24305 VDD.n802 VDD.n684 0.416
R24306 VDD.n806 VDD.n684 0.416
R24307 VDD.n807 VDD.n806 0.416
R24308 VDD.n807 VDD.n682 0.416
R24309 VDD.n811 VDD.n682 0.416
R24310 VDD.n812 VDD.n811 0.416
R24311 VDD.n812 VDD.n680 0.416
R24312 VDD.n816 VDD.n680 0.416
R24313 VDD.n817 VDD.n816 0.416
R24314 VDD.n817 VDD.n678 0.416
R24315 VDD.n821 VDD.n678 0.416
R24316 VDD.n822 VDD.n821 0.416
R24317 VDD.n824 VDD.n822 0.416
R24318 VDD.n824 VDD.n823 0.416
R24319 VDD.n823 VDD.n673 0.416
R24320 VDD.n831 VDD.n673 0.416
R24321 VDD.n834 VDD.n833 0.416
R24322 VDD.n834 VDD.n671 0.416
R24323 VDD.n839 VDD.n671 0.416
R24324 VDD.n840 VDD.n839 0.416
R24325 VDD.n841 VDD.n840 0.416
R24326 VDD.n841 VDD.n667 0.416
R24327 VDD.n847 VDD.n667 0.416
R24328 VDD.n460 VDD.n458 0.416
R24329 VDD.n464 VDD.n460 0.416
R24330 VDD.n466 VDD.n464 0.416
R24331 VDD.n468 VDD.n466 0.416
R24332 VDD.n470 VDD.n468 0.416
R24333 VDD.n474 VDD.n470 0.416
R24334 VDD.n476 VDD.n474 0.416
R24335 VDD.n478 VDD.n476 0.416
R24336 VDD.n482 VDD.n478 0.416
R24337 VDD.n484 VDD.n482 0.416
R24338 VDD.n486 VDD.n484 0.416
R24339 VDD.n490 VDD.n486 0.416
R24340 VDD.n492 VDD.n490 0.416
R24341 VDD.n494 VDD.n492 0.416
R24342 VDD.n498 VDD.n494 0.416
R24343 VDD.n500 VDD.n498 0.416
R24344 VDD.n502 VDD.n500 0.416
R24345 VDD.n504 VDD.n502 0.416
R24346 VDD.n508 VDD.n504 0.416
R24347 VDD.n510 VDD.n508 0.416
R24348 VDD.n512 VDD.n510 0.416
R24349 VDD.n516 VDD.n512 0.416
R24350 VDD.n518 VDD.n516 0.416
R24351 VDD.n520 VDD.n518 0.416
R24352 VDD.n524 VDD.n520 0.416
R24353 VDD.n526 VDD.n524 0.416
R24354 VDD.n528 VDD.n526 0.416
R24355 VDD.n532 VDD.n528 0.416
R24356 VDD.n534 VDD.n532 0.416
R24357 VDD.n536 VDD.n534 0.416
R24358 VDD.n538 VDD.n536 0.416
R24359 VDD.n542 VDD.n538 0.416
R24360 VDD.n544 VDD.n542 0.416
R24361 VDD.n546 VDD.n544 0.416
R24362 VDD.n550 VDD.n546 0.416
R24363 VDD.n552 VDD.n550 0.416
R24364 VDD.n554 VDD.n552 0.416
R24365 VDD.n558 VDD.n554 0.416
R24366 VDD.n560 VDD.n558 0.416
R24367 VDD.n562 VDD.n560 0.416
R24368 VDD.n566 VDD.n562 0.416
R24369 VDD.n568 VDD.n566 0.416
R24370 VDD.n570 VDD.n568 0.416
R24371 VDD.n572 VDD.n570 0.416
R24372 VDD.n576 VDD.n572 0.416
R24373 VDD.n578 VDD.n576 0.416
R24374 VDD.n580 VDD.n578 0.416
R24375 VDD.n584 VDD.n580 0.416
R24376 VDD.n586 VDD.n584 0.416
R24377 VDD.n588 VDD.n586 0.416
R24378 VDD.n595 VDD.n593 0.416
R24379 VDD.n597 VDD.n595 0.416
R24380 VDD.n601 VDD.n597 0.416
R24381 VDD.n603 VDD.n601 0.416
R24382 VDD.n605 VDD.n603 0.416
R24383 VDD.n607 VDD.n605 0.416
R24384 VDD.n611 VDD.n607 0.416
R24385 VDD.n613 VDD.n611 0.416
R24386 VDD.n615 VDD.n613 0.416
R24387 VDD.n619 VDD.n615 0.416
R24388 VDD.n621 VDD.n619 0.416
R24389 VDD.n624 VDD.n621 0.416
R24390 VDD.n629 VDD.n628 0.416
R24391 VDD.n628 VDD.n627 0.416
R24392 VDD.n627 VDD.n236 0.416
R24393 VDD.n637 VDD.n236 0.416
R24394 VDD.n638 VDD.n637 0.416
R24395 VDD.n639 VDD.n638 0.416
R24396 VDD.n639 VDD.n233 0.416
R24397 VDD.n645 VDD.n233 0.416
R24398 VDD.n1190 VDD.n1189 0.416
R24399 VDD.n1189 VDD.n186 0.416
R24400 VDD.n1185 VDD.n186 0.416
R24401 VDD.n1182 VDD.n190 0.416
R24402 VDD.n1178 VDD.n190 0.416
R24403 VDD.n1424 VDD.n1422 0.416
R24404 VDD.n1422 VDD.n1420 0.416
R24405 VDD.n1420 VDD.n1416 0.416
R24406 VDD.n1416 VDD.n1414 0.416
R24407 VDD.n1414 VDD.n1412 0.416
R24408 VDD.n1412 VDD.n1410 0.416
R24409 VDD.n1410 VDD.n1406 0.416
R24410 VDD.n1406 VDD.n1404 0.416
R24411 VDD.n1404 VDD.n1402 0.416
R24412 VDD.n1402 VDD.n1398 0.416
R24413 VDD.n1398 VDD.n1396 0.416
R24414 VDD.n1396 VDD.n1394 0.416
R24415 VDD.n1394 VDD.n1390 0.416
R24416 VDD.n1390 VDD.n1388 0.416
R24417 VDD.n1388 VDD.n1386 0.416
R24418 VDD.n1386 VDD.n1382 0.416
R24419 VDD.n1382 VDD.n1380 0.416
R24420 VDD.n1380 VDD.n1378 0.416
R24421 VDD.n1378 VDD.n1376 0.416
R24422 VDD.n1376 VDD.n1372 0.416
R24423 VDD.n1372 VDD.n1370 0.416
R24424 VDD.n1370 VDD.n1368 0.416
R24425 VDD.n1368 VDD.n1364 0.416
R24426 VDD.n1364 VDD.n1362 0.416
R24427 VDD.n1362 VDD.n1360 0.416
R24428 VDD.n1360 VDD.n1356 0.416
R24429 VDD.n1356 VDD.n1354 0.416
R24430 VDD.n1354 VDD.n1352 0.416
R24431 VDD.n1352 VDD.n1348 0.416
R24432 VDD.n1348 VDD.n1346 0.416
R24433 VDD.n1346 VDD.n1344 0.416
R24434 VDD.n1344 VDD.n1342 0.416
R24435 VDD.n1342 VDD.n1338 0.416
R24436 VDD.n1338 VDD.n1336 0.416
R24437 VDD.n1336 VDD.n1334 0.416
R24438 VDD.n1334 VDD.n1330 0.416
R24439 VDD.n1330 VDD.n1328 0.416
R24440 VDD.n1328 VDD.n1326 0.416
R24441 VDD.n1326 VDD.n1322 0.416
R24442 VDD.n1322 VDD.n1320 0.416
R24443 VDD.n1320 VDD.n1318 0.416
R24444 VDD.n1318 VDD.n1314 0.416
R24445 VDD.n1314 VDD.n1312 0.416
R24446 VDD.n1312 VDD.n1310 0.416
R24447 VDD.n1310 VDD.n1308 0.416
R24448 VDD.n1308 VDD.n1304 0.416
R24449 VDD.n1487 VDD.n1483 0.416
R24450 VDD.n1489 VDD.n1487 0.416
R24451 VDD.n1491 VDD.n1489 0.416
R24452 VDD.n1495 VDD.n1491 0.416
R24453 VDD.n1497 VDD.n1495 0.416
R24454 VDD.n1499 VDD.n1497 0.416
R24455 VDD.n1503 VDD.n1499 0.416
R24456 VDD.n1505 VDD.n1503 0.416
R24457 VDD.n1510 VDD.n1508 0.416
R24458 VDD.n1514 VDD.n1510 0.416
R24459 VDD.n1516 VDD.n1514 0.416
R24460 VDD.n1518 VDD.n1516 0.416
R24461 VDD.n1522 VDD.n1518 0.416
R24462 VDD.n1524 VDD.n1522 0.416
R24463 VDD.n1527 VDD.n1524 0.416
R24464 VDD.n362 VDD.n361 0.376
R24465 VDD.n346 VDD.n345 0.376
R24466 VDD.n904 VDD.n868 0.337
R24467 VDD.n589 VDD.n588 0.308
R24468 VDD.n1192 VDD.n1191 0.28
R24469 VDD.n1508 VDD.n1506 0.275
R24470 VDD.n1183 VDD.n1182 0.227
R24471 VDD.n1274 VDD.n0 0.226
R24472 VDD.n195 VDD.n194 0.226
R24473 VDD.n1561 VDD.n1560 0.226
R24474 VDD.n0  0.218
R24475  VDD.n1561 0.218
R24476 VDD.n1211 VDD.n1210 0.217
R24477 VDD.n1216 VDD.n1215 0.217
R24478 VDD.n1221 VDD.n1220 0.217
R24479 VDD.n1226 VDD.n1225 0.217
R24480 VDD.n1231 VDD.n1230 0.217
R24481 VDD.n1236 VDD.n1235 0.217
R24482 VDD.n1241 VDD.n1240 0.217
R24483 VDD.n1246 VDD.n1245 0.217
R24484 VDD.n1251 VDD.n1250 0.217
R24485 VDD.n1435 VDD.n1434 0.217
R24486 VDD.n1161 VDD.n1160 0.217
R24487 VDD.n1150 VDD.n1149 0.217
R24488 VDD.n1139 VDD.n1138 0.217
R24489 VDD.n1128 VDD.n1127 0.217
R24490 VDD.n1118 VDD.n1117 0.217
R24491 VDD.n1108 VDD.n1107 0.217
R24492 VDD.n1097 VDD.n1096 0.217
R24493 VDD.n1087 VDD.n1086 0.217
R24494 VDD.n1076 VDD.n1075 0.217
R24495 VDD.n1480 VDD.n1479 0.217
R24496 VDD.n1184 VDD.n1183 0.211
R24497 VDD.n832 VDD.n831 0.208
R24498 VDD.n833 VDD.n832 0.208
R24499 VDD.n358 VDD.n355 0.19
R24500 VDD.n193  0.174
R24501 VDD.n194  0.174
R24502 VDD.n274 VDD.n271 0.163
R24503 VDD.n1191 VDD.n1190 0.158
R24504 VDD.n436 VDD.n434 0.144
R24505 VDD.n425 VDD.n423 0.144
R24506 VDD.n414 VDD.n412 0.144
R24507 VDD.n403 VDD.n401 0.144
R24508 VDD.n392 VDD.n390 0.144
R24509 VDD.n381 VDD.n379 0.144
R24510 VDD.n370 VDD.n368 0.144
R24511 VDD.n351 VDD.n344 0.144
R24512 VDD.n340 VDD.n333 0.144
R24513 VDD.n329 VDD.n322 0.144
R24514 VDD.n318 VDD.n311 0.144
R24515 VDD.n307 VDD.n300 0.144
R24516 VDD.n296 VDD.n289 0.144
R24517 VDD.n285 VDD.n278 0.144
R24518 VDD.n1506 VDD.n1505 0.141
R24519 VDD.n1561 VDD 0.137
R24520 VDD.n194  0.137
R24521 VDD.n0  0.11
R24522 VDD.n193  0.11
R24523 VDD.n593 VDD.n589 0.108
R24524 VDD.n897 VDD.n868 0.079
R24525 VDD.n1049 VDD.n1044 0.077
R24526 VDD.n1017 VDD.n1012 0.077
R24527 VDD.n986 VDD.n981 0.077
R24528 VDD.n954 VDD.n949 0.077
R24529 VDD.n917 VDD.n912 0.077
R24530 VDD.n860 VDD.n855 0.077
R24531 VDD.n659 VDD.n654 0.077
R24532 VDD.n213 VDD.n208 0.077
R24533 VDD.n202 VDD.n197 0.077
R24534 VDD.n1467 VDD.n1462 0.077
R24535 VDD.n1272 VDD.n1271 0.077
R24536 VDD.n1555 VDD.n1554 0.076
R24537 VDD.n11 VDD.n10 0.076
R24538 VDD.n32 VDD.n31 0.076
R24539 VDD.n53 VDD.n52 0.076
R24540 VDD.n74 VDD.n73 0.076
R24541 VDD.n95 VDD.n94 0.076
R24542 VDD.n116 VDD.n115 0.076
R24543 VDD.n137 VDD.n136 0.076
R24544 VDD.n158 VDD.n157 0.076
R24545 VDD.n177 VDD.n172 0.076
R24546 VDD.n1284 VDD.n1283 0.076
R24547 VDD.n1068 VDD.n1056 0.074
R24548 VDD.n1067 VDD.n1057 0.074
R24549 VDD.n1037 VDD.n1025 0.074
R24550 VDD.n1036 VDD.n1026 0.074
R24551 VDD.n1005 VDD.n993 0.074
R24552 VDD.n1004 VDD.n994 0.074
R24553 VDD.n974 VDD.n962 0.074
R24554 VDD.n973 VDD.n963 0.074
R24555 VDD.n942 VDD.n925 0.074
R24556 VDD.n936 VDD.n926 0.074
R24557 VDD.n905 VDD.n867 0.074
R24558 VDD.n884 VDD.n874 0.074
R24559 VDD.n848 VDD.n666 0.074
R24560 VDD.n726 VDD.n716 0.074
R24561 VDD.n647 VDD.n220 0.074
R24562 VDD.n454 VDD.n444 0.074
R24563 VDD.n1177 VDD.n1176 0.074
R24564 VDD.n1193 VDD.n184 0.074
R24565 VDD.n1450 VDD.n1449 0.074
R24566 VDD.n1529 VDD.n1528 0.074
R24567 VDD.n368 VDD.n360 0.043
R24568 VDD.n353 VDD.n351 0.043
R24569 VDD.n1447 VDD.n1446 0.042
R24570 VDD.n1428 VDD.n1427 0.042
R24571 VDD.n1445 VDD.n1444 0.041
R24572 VDD.n1429 VDD.n1301 0.041
R24573 VDD.n438 VDD.n436 0.04
R24574 VDD.n278 VDD.n276 0.04
R24575 VDD.n379 VDD.n372 0.038
R24576 VDD.n342 VDD.n340 0.038
R24577 VDD.n1444 VDD.n1443 0.036
R24578 VDD.n1301 VDD.n1300 0.036
R24579 VDD.n1448 VDD.n1447 0.036
R24580 VDD.n1427 VDD.n1426 0.036
R24581 VDD.n427 VDD.n425 0.035
R24582 VDD.n289 VDD.n287 0.035
R24583 VDD.n390 VDD.n383 0.032
R24584 VDD.n331 VDD.n329 0.032
R24585 VDD.n416 VDD.n414 0.029
R24586 VDD.n300 VDD.n298 0.029
R24587 VDD.n401 VDD.n394 0.027
R24588 VDD.n320 VDD.n318 0.027
R24589 VDD.n405 VDD.n403 0.024
R24590 VDD.n311 VDD.n309 0.024
R24591 VDD.n1204 VDD.n1203 0.024
R24592 VDD.n1206 VDD.n1205 0.024
R24593 VDD.n1537 VDD.n1534 0.024
R24594 VDD.n1475 VDD.n1474 0.024
R24595 VDD.n1473 VDD.n1472 0.024
R24596 VDD.n1273 VDD.n1272 0.023
R24597 VDD.n1064 VDD.n1063 0.021
R24598 VDD.n1033 VDD.n1032 0.021
R24599 VDD.n1001 VDD.n1000 0.021
R24600 VDD.n970 VDD.n969 0.021
R24601 VDD.n933 VDD.n932 0.021
R24602 VDD.n881 VDD.n880 0.021
R24603 VDD.n723 VDD.n722 0.021
R24604 VDD.n451 VDD.n450 0.021
R24605 VDD.n13 VDD.n5 0.021
R24606 VDD.n4 VDD.n2 0.021
R24607 VDD.n1064 VDD.n1062 0.021
R24608 VDD.n34 VDD.n26 0.021
R24609 VDD.n25 VDD.n23 0.021
R24610 VDD.n1033 VDD.n1031 0.021
R24611 VDD.n55 VDD.n47 0.021
R24612 VDD.n46 VDD.n44 0.021
R24613 VDD.n1001 VDD.n999 0.021
R24614 VDD.n76 VDD.n68 0.021
R24615 VDD.n67 VDD.n65 0.021
R24616 VDD.n970 VDD.n968 0.021
R24617 VDD.n97 VDD.n89 0.021
R24618 VDD.n88 VDD.n86 0.021
R24619 VDD.n933 VDD.n931 0.021
R24620 VDD.n118 VDD.n110 0.021
R24621 VDD.n109 VDD.n107 0.021
R24622 VDD.n881 VDD.n879 0.021
R24623 VDD.n139 VDD.n131 0.021
R24624 VDD.n130 VDD.n128 0.021
R24625 VDD.n723 VDD.n721 0.021
R24626 VDD.n160 VDD.n152 0.021
R24627 VDD.n151 VDD.n149 0.021
R24628 VDD.n451 VDD.n449 0.021
R24629 VDD.n412 VDD.n405 0.021
R24630 VDD.n309 VDD.n307 0.021
R24631 VDD.n176 VDD.n175 0.021
R24632 VDD.n1080 VDD.n1079 0.021
R24633 VDD.n1101 VDD.n1100 0.021
R24634 VDD.n1132 VDD.n1131 0.021
R24635 VDD.n1143 VDD.n1142 0.021
R24636 VDD.n1154 VDD.n1153 0.021
R24637 VDD.n1165 VDD.n1164 0.021
R24638 VDD.n1022 VDD.n1021 0.021
R24639 VDD.n959 VDD.n958 0.021
R24640 VDD.n922 VDD.n921 0.021
R24641 VDD.n1061 VDD.n1060 0.021
R24642 VDD.n1030 VDD.n1029 0.021
R24643 VDD.n998 VDD.n997 0.021
R24644 VDD.n967 VDD.n966 0.021
R24645 VDD.n930 VDD.n929 0.021
R24646 VDD.n878 VDD.n877 0.021
R24647 VDD.n720 VDD.n719 0.021
R24648 VDD.n448 VDD.n447 0.021
R24649 VDD.n1207 VDD.n181 0.019
R24650 VDD.n1476 VDD.n1459 0.019
R24651 VDD.n394 VDD.n392 0.019
R24652 VDD.n322 VDD.n320 0.019
R24653 VDD.n1072 VDD.n1071 0.018
R24654 VDD.n1041 VDD.n1040 0.018
R24655 VDD.n1009 VDD.n1008 0.018
R24656 VDD.n978 VDD.n977 0.018
R24657 VDD.n946 VDD.n945 0.018
R24658 VDD.n909 VDD.n908 0.018
R24659 VDD.n852 VDD.n851 0.018
R24660 VDD.n651 VDD.n650 0.018
R24661 VDD.n1174 VDD.n1173 0.018
R24662 VDD.n1197 VDD.n1196 0.018
R24663 VDD.n1454 VDD.n1453 0.018
R24664 VDD.n1466 VDD.n1465 0.018
R24665 VDD.n1533 VDD.n1532 0.018
R24666 VDD.n1431 VDD.n1430 0.018
R24667 VDD.n1295 VDD.n1294 0.018
R24668 VDD.n1290 VDD.n1289 0.018
R24669 VDD.n1285 VDD.n1284 0.018
R24670 VDD.n14 VDD.n13 0.017
R24671 VDD.n20 VDD.n19 0.017
R24672 VDD.n22 VDD.n21 0.017
R24673 VDD.n35 VDD.n34 0.017
R24674 VDD.n41 VDD.n40 0.017
R24675 VDD.n43 VDD.n42 0.017
R24676 VDD.n56 VDD.n55 0.017
R24677 VDD.n62 VDD.n61 0.017
R24678 VDD.n64 VDD.n63 0.017
R24679 VDD.n77 VDD.n76 0.017
R24680 VDD.n83 VDD.n82 0.017
R24681 VDD.n85 VDD.n84 0.017
R24682 VDD.n98 VDD.n97 0.017
R24683 VDD.n104 VDD.n103 0.017
R24684 VDD.n106 VDD.n105 0.017
R24685 VDD.n119 VDD.n118 0.017
R24686 VDD.n125 VDD.n124 0.017
R24687 VDD.n127 VDD.n126 0.017
R24688 VDD.n140 VDD.n139 0.017
R24689 VDD.n146 VDD.n145 0.017
R24690 VDD.n148 VDD.n147 0.017
R24691 VDD.n161 VDD.n160 0.017
R24692 VDD.n167 VDD.n166 0.017
R24693 VDD.n169 VDD.n168 0.017
R24694 VDD.n1285 VDD.n1278 0.016
R24695 VDD.n1290 VDD.n1288 0.016
R24696 VDD.n1295 VDD.n1293 0.016
R24697 VDD.n1431 VDD.n1429 0.016
R24698 VDD.n423 VDD.n416 0.016
R24699 VDD.n298 VDD.n296 0.016
R24700 VDD.n14 VDD.n4 0.016
R24701 VDD.n20 VDD.n17 0.016
R24702 VDD.n1064 VDD.n22 0.016
R24703 VDD.n35 VDD.n25 0.016
R24704 VDD.n41 VDD.n38 0.016
R24705 VDD.n1033 VDD.n43 0.016
R24706 VDD.n56 VDD.n46 0.016
R24707 VDD.n62 VDD.n59 0.016
R24708 VDD.n1001 VDD.n64 0.016
R24709 VDD.n77 VDD.n67 0.016
R24710 VDD.n83 VDD.n80 0.016
R24711 VDD.n970 VDD.n85 0.016
R24712 VDD.n98 VDD.n88 0.016
R24713 VDD.n104 VDD.n101 0.016
R24714 VDD.n933 VDD.n106 0.016
R24715 VDD.n119 VDD.n109 0.016
R24716 VDD.n125 VDD.n122 0.016
R24717 VDD.n881 VDD.n127 0.016
R24718 VDD.n140 VDD.n130 0.016
R24719 VDD.n146 VDD.n143 0.016
R24720 VDD.n723 VDD.n148 0.016
R24721 VDD.n161 VDD.n151 0.016
R24722 VDD.n167 VDD.n164 0.016
R24723 VDD.n451 VDD.n169 0.016
R24724 VDD.n1284 VDD.n1282 0.015
R24725 VDD.n1278 VDD.n1276 0.015
R24726 VDD.n1288 VDD.n1286 0.015
R24727 VDD.n1293 VDD.n1291 0.015
R24728 VDD.n1429 VDD.n1299 0.015
R24729 VDD.n1049 VDD.n1048 0.015
R24730 VDD.n11 VDD.n9 0.015
R24731 VDD.n12 VDD.n11 0.015
R24732 VDD.n13 VDD.n12 0.015
R24733 VDD.n4 VDD.n3 0.015
R24734 VDD.n17 VDD.n15 0.015
R24735 VDD.n1065 VDD.n1064 0.015
R24736 VDD.n1066 VDD.n1065 0.015
R24737 VDD.n1017 VDD.n1016 0.015
R24738 VDD.n32 VDD.n30 0.015
R24739 VDD.n33 VDD.n32 0.015
R24740 VDD.n34 VDD.n33 0.015
R24741 VDD.n25 VDD.n24 0.015
R24742 VDD.n38 VDD.n36 0.015
R24743 VDD.n1034 VDD.n1033 0.015
R24744 VDD.n1035 VDD.n1034 0.015
R24745 VDD.n986 VDD.n985 0.015
R24746 VDD.n53 VDD.n51 0.015
R24747 VDD.n54 VDD.n53 0.015
R24748 VDD.n55 VDD.n54 0.015
R24749 VDD.n46 VDD.n45 0.015
R24750 VDD.n59 VDD.n57 0.015
R24751 VDD.n1002 VDD.n1001 0.015
R24752 VDD.n1003 VDD.n1002 0.015
R24753 VDD.n954 VDD.n953 0.015
R24754 VDD.n74 VDD.n72 0.015
R24755 VDD.n75 VDD.n74 0.015
R24756 VDD.n76 VDD.n75 0.015
R24757 VDD.n67 VDD.n66 0.015
R24758 VDD.n80 VDD.n78 0.015
R24759 VDD.n971 VDD.n970 0.015
R24760 VDD.n972 VDD.n971 0.015
R24761 VDD.n917 VDD.n916 0.015
R24762 VDD.n95 VDD.n93 0.015
R24763 VDD.n96 VDD.n95 0.015
R24764 VDD.n97 VDD.n96 0.015
R24765 VDD.n88 VDD.n87 0.015
R24766 VDD.n101 VDD.n99 0.015
R24767 VDD.n934 VDD.n933 0.015
R24768 VDD.n935 VDD.n934 0.015
R24769 VDD.n860 VDD.n859 0.015
R24770 VDD.n116 VDD.n114 0.015
R24771 VDD.n117 VDD.n116 0.015
R24772 VDD.n118 VDD.n117 0.015
R24773 VDD.n109 VDD.n108 0.015
R24774 VDD.n122 VDD.n120 0.015
R24775 VDD.n882 VDD.n881 0.015
R24776 VDD.n883 VDD.n882 0.015
R24777 VDD.n659 VDD.n658 0.015
R24778 VDD.n137 VDD.n135 0.015
R24779 VDD.n138 VDD.n137 0.015
R24780 VDD.n139 VDD.n138 0.015
R24781 VDD.n130 VDD.n129 0.015
R24782 VDD.n143 VDD.n141 0.015
R24783 VDD.n724 VDD.n723 0.015
R24784 VDD.n725 VDD.n724 0.015
R24785 VDD.n213 VDD.n212 0.015
R24786 VDD.n158 VDD.n156 0.015
R24787 VDD.n159 VDD.n158 0.015
R24788 VDD.n160 VDD.n159 0.015
R24789 VDD.n151 VDD.n150 0.015
R24790 VDD.n164 VDD.n162 0.015
R24791 VDD.n452 VDD.n451 0.015
R24792 VDD.n453 VDD.n452 0.015
R24793 VDD.n202 VDD.n201 0.015
R24794 VDD.n1272 VDD.n1270 0.015
R24795 VDD.n1445 VDD.n1442 0.015
R24796 VDD.n1556 VDD.n1553 0.015
R24797 VDD.n1074 VDD.n1073 0.014
R24798 VDD.n1043 VDD.n1042 0.014
R24799 VDD.n1011 VDD.n1010 0.014
R24800 VDD.n980 VDD.n979 0.014
R24801 VDD.n948 VDD.n947 0.014
R24802 VDD.n911 VDD.n910 0.014
R24803 VDD.n854 VDD.n853 0.014
R24804 VDD.n653 VDD.n652 0.014
R24805 VDD.n1175 VDD.n1170 0.014
R24806 VDD.n1207 VDD.n1206 0.013
R24807 VDD.n1476 VDD.n1475 0.013
R24808 VDD.n383 VDD.n381 0.013
R24809 VDD.n333 VDD.n331 0.013
R24810 VDD.n1282 VDD.n1281 0.013
R24811 VDD.n1299 VDD.n1298 0.013
R24812 VDD.n1048 VDD.n1047 0.013
R24813 VDD.n9 VDD.n8 0.013
R24814 VDD.n1016 VDD.n1015 0.013
R24815 VDD.n30 VDD.n29 0.013
R24816 VDD.n985 VDD.n984 0.013
R24817 VDD.n51 VDD.n50 0.013
R24818 VDD.n953 VDD.n952 0.013
R24819 VDD.n72 VDD.n71 0.013
R24820 VDD.n916 VDD.n915 0.013
R24821 VDD.n93 VDD.n92 0.013
R24822 VDD.n859 VDD.n858 0.013
R24823 VDD.n114 VDD.n113 0.013
R24824 VDD.n658 VDD.n657 0.013
R24825 VDD.n135 VDD.n134 0.013
R24826 VDD.n212 VDD.n211 0.013
R24827 VDD.n156 VDD.n155 0.013
R24828 VDD.n201 VDD.n200 0.013
R24829 VDD.n1270 VDD.n1269 0.013
R24830 VDD.n1442 VDD.n1441 0.013
R24831 VDD.n1553 VDD.n1552 0.013
R24832 VDD.n178 VDD.n177 0.012
R24833 VDD.n180 VDD.n179 0.012
R24834 VDD.n1202 VDD.n1201 0.012
R24835 VDD.n1456 VDD.n1455 0.012
R24836 VDD.n1471 VDD.n1470 0.012
R24837 VDD.n1073 VDD.n1072 0.01
R24838 VDD.n1042 VDD.n1041 0.01
R24839 VDD.n1010 VDD.n1009 0.01
R24840 VDD.n979 VDD.n978 0.01
R24841 VDD.n947 VDD.n946 0.01
R24842 VDD.n910 VDD.n909 0.01
R24843 VDD.n853 VDD.n852 0.01
R24844 VDD.n652 VDD.n651 0.01
R24845 VDD.n1175 VDD.n1174 0.01
R24846 VDD.n1198 VDD.n1197 0.01
R24847 VDD.n1455 VDD.n1454 0.01
R24848 VDD.n1534 VDD.n1533 0.01
R24849 VDD.n1467 VDD.n1466 0.01
R24850 VDD.n434 VDD.n427 0.01
R24851 VDD.n287 VDD.n285 0.01
R24852 VDD.n1199 VDD.n1198 0.01
R24853 VDD.n1459 VDD.n1458 0.01
R24854 VDD.n1468 VDD.n1467 0.01
R24855 VDD.n1200 VDD.n1199 0.009
R24856 VDD.n1458 VDD.n1457 0.009
R24857 VDD.n1469 VDD.n1468 0.009
R24858 VDD.n453 VDD.n448 0.008
R24859 VDD.n725 VDD.n720 0.008
R24860 VDD.n883 VDD.n878 0.008
R24861 VDD.n935 VDD.n930 0.008
R24862 VDD.n972 VDD.n967 0.008
R24863 VDD.n1003 VDD.n998 0.008
R24864 VDD.n1035 VDD.n1030 0.008
R24865 VDD.n1066 VDD.n1061 0.008
R24866 VDD.n1081 VDD.n1080 0.008
R24867 VDD.n1091 VDD.n1090 0.008
R24868 VDD.n1102 VDD.n1101 0.008
R24869 VDD.n1112 VDD.n1111 0.008
R24870 VDD.n1122 VDD.n1121 0.008
R24871 VDD.n1133 VDD.n1132 0.008
R24872 VDD.n1144 VDD.n1143 0.008
R24873 VDD.n1155 VDD.n1154 0.008
R24874 VDD.n1166 VDD.n1165 0.008
R24875 VDD.n1205 VDD.n1204 0.008
R24876 VDD.n1203 VDD.n1202 0.008
R24877 VDD.n1474 VDD.n1473 0.008
R24878 VDD.n1472 VDD.n1471 0.008
R24879 VDD.n1537 VDD.n1536 0.008
R24880 VDD.n1539 VDD.n1538 0.008
R24881 VDD.n1542 VDD.n1541 0.008
R24882 VDD.n1544 VDD.n1543 0.008
R24883 VDD.n1547 VDD.n1546 0.008
R24884 VDD.n1549 VDD.n1548 0.008
R24885 VDD.n1557 VDD.n1556 0.008
R24886 VDD.n372 VDD.n370 0.008
R24887 VDD.n344 VDD.n342 0.008
R24888 VDD.n177 VDD.n176 0.008
R24889 VDD.n1445 VDD.n1438 0.008
R24890 VDD.n1254 VDD.n1253 0.008
R24891 VDD.n1257 VDD.n1256 0.008
R24892 VDD.n1259 VDD.n1258 0.008
R24893 VDD.n1262 VDD.n1261 0.008
R24894 VDD.n1264 VDD.n1263 0.008
R24895 VDD.n1273 VDD.n1266 0.008
R24896 VDD.n179 VDD.n178 0.007
R24897 VDD.n181 VDD.n180 0.007
R24898 VDD.n1201 VDD.n1200 0.007
R24899 VDD.n1470 VDD.n1469 0.007
R24900 VDD.n1457 VDD.n1456 0.007
R24901 VDD.n646 VDD.n645 0.006
R24902 VDD.n1074 VDD.n1055 0.005
R24903 VDD.n1083 VDD.n1082 0.005
R24904 VDD.n1054 VDD.n1053 0.005
R24905 VDD.n1052 VDD.n1051 0.005
R24906 VDD.n1078 VDD.n1077 0.005
R24907 VDD.n1050 VDD.n1049 0.005
R24908 VDD.n1043 VDD.n1024 0.005
R24909 VDD.n1093 VDD.n1092 0.005
R24910 VDD.n1023 VDD.n1022 0.005
R24911 VDD.n1020 VDD.n1019 0.005
R24912 VDD.n1089 VDD.n1088 0.005
R24913 VDD.n1018 VDD.n1017 0.005
R24914 VDD.n1011 VDD.n992 0.005
R24915 VDD.n1104 VDD.n1103 0.005
R24916 VDD.n991 VDD.n990 0.005
R24917 VDD.n989 VDD.n988 0.005
R24918 VDD.n1099 VDD.n1098 0.005
R24919 VDD.n987 VDD.n986 0.005
R24920 VDD.n980 VDD.n961 0.005
R24921 VDD.n1114 VDD.n1113 0.005
R24922 VDD.n960 VDD.n959 0.005
R24923 VDD.n957 VDD.n956 0.005
R24924 VDD.n1110 VDD.n1109 0.005
R24925 VDD.n955 VDD.n954 0.005
R24926 VDD.n948 VDD.n924 0.005
R24927 VDD.n1124 VDD.n1123 0.005
R24928 VDD.n923 VDD.n922 0.005
R24929 VDD.n920 VDD.n919 0.005
R24930 VDD.n1120 VDD.n1119 0.005
R24931 VDD.n918 VDD.n917 0.005
R24932 VDD.n911 VDD.n866 0.005
R24933 VDD.n1135 VDD.n1134 0.005
R24934 VDD.n865 VDD.n864 0.005
R24935 VDD.n863 VDD.n862 0.005
R24936 VDD.n1130 VDD.n1129 0.005
R24937 VDD.n861 VDD.n860 0.005
R24938 VDD.n854 VDD.n665 0.005
R24939 VDD.n1146 VDD.n1145 0.005
R24940 VDD.n664 VDD.n663 0.005
R24941 VDD.n662 VDD.n661 0.005
R24942 VDD.n1141 VDD.n1140 0.005
R24943 VDD.n660 VDD.n659 0.005
R24944 VDD.n653 VDD.n219 0.005
R24945 VDD.n1157 VDD.n1156 0.005
R24946 VDD.n218 VDD.n217 0.005
R24947 VDD.n216 VDD.n215 0.005
R24948 VDD.n1152 VDD.n1151 0.005
R24949 VDD.n214 VDD.n213 0.005
R24950 VDD.n1170 VDD.n192 0.005
R24951 VDD.n1168 VDD.n1167 0.005
R24952 VDD.n207 VDD.n206 0.005
R24953 VDD.n205 VDD.n204 0.005
R24954 VDD.n1163 VDD.n1162 0.005
R24955 VDD.n203 VDD.n202 0.005
R24956 VDD.n441 VDD.n438 0.005
R24957 VDD.n276 VDD.n274 0.005
R24958 VDD.n174 VDD.n173 0.005
R24959 VDD.n1297 VDD.n1296 0.005
R24960 VDD.n1059 VDD.n1058 0.005
R24961 VDD.n1028 VDD.n1027 0.005
R24962 VDD.n996 VDD.n995 0.005
R24963 VDD.n965 VDD.n964 0.005
R24964 VDD.n928 VDD.n927 0.005
R24965 VDD.n876 VDD.n875 0.005
R24966 VDD.n718 VDD.n717 0.005
R24967 VDD.n446 VDD.n445 0.005
R24968 VDD.n1268 VDD.n1267 0.005
R24969 VDD.n1452 VDD.n1451 0.005
R24970 VDD.n1531 VDD.n1530 0.005
R24971 VDD.n1073 VDD.n1068 0.003
R24972 VDD.n1067 VDD.n1066 0.003
R24973 VDD.n1042 VDD.n1037 0.003
R24974 VDD.n1036 VDD.n1035 0.003
R24975 VDD.n1010 VDD.n1005 0.003
R24976 VDD.n1004 VDD.n1003 0.003
R24977 VDD.n979 VDD.n974 0.003
R24978 VDD.n973 VDD.n972 0.003
R24979 VDD.n947 VDD.n942 0.003
R24980 VDD.n936 VDD.n935 0.003
R24981 VDD.n910 VDD.n905 0.003
R24982 VDD.n884 VDD.n883 0.003
R24983 VDD.n853 VDD.n848 0.003
R24984 VDD.n726 VDD.n725 0.003
R24985 VDD.n652 VDD.n647 0.003
R24986 VDD.n454 VDD.n453 0.003
R24987 VDD.n1177 VDD.n1175 0.003
R24988 VDD.n1198 VDD.n1193 0.003
R24989 VDD.n1455 VDD.n1450 0.003
R24990 VDD.n1534 VDD.n1529 0.003
R24991 VDD.n1280 VDD.n1279 0.003
R24992 VDD.n1195 VDD.n1194 0.002
R24993 VDD.n1464 VDD.n1463 0.002
R24994 VDD.n1046 VDD.n1045 0.002
R24995 VDD.n1014 VDD.n1013 0.002
R24996 VDD.n983 VDD.n982 0.002
R24997 VDD.n951 VDD.n950 0.002
R24998 VDD.n914 VDD.n913 0.002
R24999 VDD.n857 VDD.n856 0.002
R25000 VDD.n656 VDD.n655 0.002
R25001 VDD.n210 VDD.n209 0.002
R25002 VDD.n199 VDD.n198 0.002
R25003 VDD.n7 VDD.n6 0.002
R25004 VDD.n28 VDD.n27 0.002
R25005 VDD.n49 VDD.n48 0.002
R25006 VDD.n70 VDD.n69 0.002
R25007 VDD.n91 VDD.n90 0.002
R25008 VDD.n112 VDD.n111 0.002
R25009 VDD.n133 VDD.n132 0.002
R25010 VDD.n154 VDD.n153 0.002
R25011 VDD.n1070 VDD.n1069 0.002
R25012 VDD.n1039 VDD.n1038 0.002
R25013 VDD.n1007 VDD.n1006 0.002
R25014 VDD.n976 VDD.n975 0.002
R25015 VDD.n944 VDD.n943 0.002
R25016 VDD.n907 VDD.n906 0.002
R25017 VDD.n850 VDD.n849 0.002
R25018 VDD.n649 VDD.n648 0.002
R25019 VDD.n1172 VDD.n1171 0.002
R25020 VDD.n1551 VDD.n1550 0.002
R25021 VDD.n1440 VDD.n1439 0.002
R25022 VDD.n360 VDD.n358 0.002
R25023 VDD.n355 VDD.n353 0.002
R25024 VDD.n1212 VDD.n1211 0.001
R25025 VDD.n1215 VDD.n1214 0.001
R25026 VDD.n1217 VDD.n1216 0.001
R25027 VDD.n1220 VDD.n1219 0.001
R25028 VDD.n1222 VDD.n1221 0.001
R25029 VDD.n1225 VDD.n1224 0.001
R25030 VDD.n1227 VDD.n1226 0.001
R25031 VDD.n1230 VDD.n1229 0.001
R25032 VDD.n1232 VDD.n1231 0.001
R25033 VDD.n1235 VDD.n1234 0.001
R25034 VDD.n1237 VDD.n1236 0.001
R25035 VDD.n1240 VDD.n1239 0.001
R25036 VDD.n1242 VDD.n1241 0.001
R25037 VDD.n1245 VDD.n1244 0.001
R25038 VDD.n1247 VDD.n1246 0.001
R25039 VDD.n1250 VDD.n1249 0.001
R25040 VDD.n1436 VDD.n1435 0.001
R25041 VDD.n1434 VDD.n1433 0.001
R25042 VDD.n1210 VDD.n1209 0.001
R25043 VDD.n1252 VDD.n1251 0.001
R25044 VDD.n1479 VDD.n1478 0.001
R25045 VDD.n1560 VDD.n1559 0.001
R25046 VDD.n1281 VDD.n1280 0.001
R25047 VDD.n1298 VDD.n1297 0.001
R25048 VDD.n1071 VDD.n1070 0.001
R25049 VDD.n1047 VDD.n1046 0.001
R25050 VDD.n8 VDD.n7 0.001
R25051 VDD.n1060 VDD.n1059 0.001
R25052 VDD.n1040 VDD.n1039 0.001
R25053 VDD.n1015 VDD.n1014 0.001
R25054 VDD.n29 VDD.n28 0.001
R25055 VDD.n1029 VDD.n1028 0.001
R25056 VDD.n1008 VDD.n1007 0.001
R25057 VDD.n984 VDD.n983 0.001
R25058 VDD.n50 VDD.n49 0.001
R25059 VDD.n997 VDD.n996 0.001
R25060 VDD.n977 VDD.n976 0.001
R25061 VDD.n952 VDD.n951 0.001
R25062 VDD.n71 VDD.n70 0.001
R25063 VDD.n966 VDD.n965 0.001
R25064 VDD.n945 VDD.n944 0.001
R25065 VDD.n915 VDD.n914 0.001
R25066 VDD.n92 VDD.n91 0.001
R25067 VDD.n929 VDD.n928 0.001
R25068 VDD.n908 VDD.n907 0.001
R25069 VDD.n858 VDD.n857 0.001
R25070 VDD.n113 VDD.n112 0.001
R25071 VDD.n877 VDD.n876 0.001
R25072 VDD.n851 VDD.n850 0.001
R25073 VDD.n657 VDD.n656 0.001
R25074 VDD.n134 VDD.n133 0.001
R25075 VDD.n719 VDD.n718 0.001
R25076 VDD.n650 VDD.n649 0.001
R25077 VDD.n211 VDD.n210 0.001
R25078 VDD.n155 VDD.n154 0.001
R25079 VDD.n447 VDD.n446 0.001
R25080 VDD.n1173 VDD.n1172 0.001
R25081 VDD.n200 VDD.n199 0.001
R25082 VDD.n175 VDD.n174 0.001
R25083 VDD.n1196 VDD.n1195 0.001
R25084 VDD.n1269 VDD.n1268 0.001
R25085 VDD.n1441 VDD.n1440 0.001
R25086 VDD.n1453 VDD.n1452 0.001
R25087 VDD.n1465 VDD.n1464 0.001
R25088 VDD.n1532 VDD.n1531 0.001
R25089 VDD.n1552 VDD.n1551 0.001
R25090 VDD.n1169 VDD.n1161 0.001
R25091 VDD.n1158 VDD.n1150 0.001
R25092 VDD.n1147 VDD.n1139 0.001
R25093 VDD.n1136 VDD.n1128 0.001
R25094 VDD.n1125 VDD.n1118 0.001
R25095 VDD.n1115 VDD.n1108 0.001
R25096 VDD.n1105 VDD.n1097 0.001
R25097 VDD.n1094 VDD.n1087 0.001
R25098 VDD.n1084 VDD.n1076 0.001
R25099 VDD.n1208 VDD.n171 0.001
R25100 VDD.n1275 VDD.n1274 0.001
R25101 VDD.n171 VDD.n170 0.001
R25102 VDD.n1432 VDD.n1275 0.001
R25103 VDD.n1169 VDD.n196 0.001
R25104 VDD.n1159 VDD.n1158 0.001
R25105 VDD.n1148 VDD.n1147 0.001
R25106 VDD.n1137 VDD.n1136 0.001
R25107 VDD.n1126 VDD.n1125 0.001
R25108 VDD.n1116 VDD.n1115 0.001
R25109 VDD.n1106 VDD.n1105 0.001
R25110 VDD.n1095 VDD.n1094 0.001
R25111 VDD.n1085 VDD.n1084 0.001
R25112 VDD.n1477 VDD.n1 0.001
R25113 VDD.n1558 VDD.n1481 0.001
R25114 VDD.n1481 VDD.n1480 0.001
R25115 VDD.n1075 VDD.n1 0.001
R25116 VDD.n1086 VDD.n1085 0.001
R25117 VDD.n1096 VDD.n1095 0.001
R25118 VDD.n1107 VDD.n1106 0.001
R25119 VDD.n1117 VDD.n1116 0.001
R25120 VDD.n1127 VDD.n1126 0.001
R25121 VDD.n1138 VDD.n1137 0.001
R25122 VDD.n1149 VDD.n1148 0.001
R25123 VDD.n1160 VDD.n1159 0.001
R25124 VDD.n196 VDD.n195 0.001
R25125 VDD.n1209 VDD.n1208 0.001
R25126 VDD.n1437 VDD.n1252 0.001
R25127 VDD.n1213 VDD.n1212 0.001
R25128 VDD.n1214 VDD.n1213 0.001
R25129 VDD.n1218 VDD.n1217 0.001
R25130 VDD.n1219 VDD.n1218 0.001
R25131 VDD.n1223 VDD.n1222 0.001
R25132 VDD.n1224 VDD.n1223 0.001
R25133 VDD.n1228 VDD.n1227 0.001
R25134 VDD.n1229 VDD.n1228 0.001
R25135 VDD.n1233 VDD.n1232 0.001
R25136 VDD.n1234 VDD.n1233 0.001
R25137 VDD.n1238 VDD.n1237 0.001
R25138 VDD.n1239 VDD.n1238 0.001
R25139 VDD.n1243 VDD.n1242 0.001
R25140 VDD.n1244 VDD.n1243 0.001
R25141 VDD.n1248 VDD.n1247 0.001
R25142 VDD.n1249 VDD.n1248 0.001
R25143 VDD.n1433 VDD.n1432 0.001
R25144 VDD.n1437 VDD.n1436 0.001
R25145 VDD.n1559 VDD.n1558 0.001
R25146 VDD.n1478 VDD.n1477 0.001
R25147 VDD.n1266 VDD.n1265 0.001
R25148 VDD.n1256 VDD.n1255 0.001
R25149 VDD.n1278 VDD.n1277 0.001
R25150 VDD.n1293 VDD.n1292 0.001
R25151 VDD.n19 VDD.n18 0.001
R25152 VDD.n17 VDD.n16 0.001
R25153 VDD.n40 VDD.n39 0.001
R25154 VDD.n38 VDD.n37 0.001
R25155 VDD.n61 VDD.n60 0.001
R25156 VDD.n59 VDD.n58 0.001
R25157 VDD.n82 VDD.n81 0.001
R25158 VDD.n80 VDD.n79 0.001
R25159 VDD.n103 VDD.n102 0.001
R25160 VDD.n101 VDD.n100 0.001
R25161 VDD.n124 VDD.n123 0.001
R25162 VDD.n122 VDD.n121 0.001
R25163 VDD.n145 VDD.n144 0.001
R25164 VDD.n143 VDD.n142 0.001
R25165 VDD.n166 VDD.n165 0.001
R25166 VDD.n164 VDD.n163 0.001
R25167 VDD.n1204 VDD.n183 0.001
R25168 VDD.n1206 VDD.n182 0.001
R25169 VDD.n1475 VDD.n1460 0.001
R25170 VDD.n1473 VDD.n1461 0.001
R25171 VDD.n1536 VDD.n1535 0.001
R25172 VDD.n1546 VDD.n1545 0.001
R25173 VDD.n1261 VDD.n1260 0.001
R25174 VDD.n1541 VDD.n1540 0.001
R25175 VDD.n1288 VDD.n1287 0.001
R25176 VDD.n1556 VDD.n1555 0.001
R25177 VDD.n1446 VDD.n1445 0.001
R25178 VDD.n1429 VDD.n1428 0.001
R25179 vb.n178 vb.n177 3161.95
R25180 vb.n0 vb.t7 244.947
R25181 vb.n192 vb.t1 218.92
R25182 vb.n189 vb.t8 218.92
R25183 vb.n3 vb.t6 218.92
R25184 vb.n186 vb.t5 218.92
R25185 vb.n2 vb.t3 218.92
R25186 vb.n183 vb.t4 218.92
R25187 vb.n1 vb.t2 218.92
R25188 vb.n179 vb.t0 218.919
R25189 vb.n100 vb.n97 176.62
R25190 vb.n184 vb.n183 105.076
R25191 vb.n198 vb.n197 85.333
R25192 vb.n197 vb.n196 85.333
R25193 vb.n196 vb.n195 85.333
R25194 vb.n195 vb.n194 85.333
R25195 vb.n194 vb.n191 85.333
R25196 vb.n191 vb.n188 85.333
R25197 vb.n188 vb.n185 85.333
R25198 vb.n185 vb.n182 85.333
R25199 vb.n182 vb.n180 85.333
R25200 vb.n180 vb.n179 78.892
R25201 vb.n187 vb.n186 78.084
R25202 vb.n198 vb.n0 76
R25203 vb.n197 vb.n1 76
R25204 vb.n196 vb.n2 76
R25205 vb.n195 vb.n3 76
R25206 vb.n194 vb.n193 76
R25207 vb.n191 vb.n190 76
R25208 vb.n188 vb.n187 76
R25209 vb.n185 vb.n184 76
R25210 vb.n182 vb.n181 76
R25211 vb.n4 vb 70.67
R25212 vb vb.n198 68.266
R25213 vb.n5 vb 60.649
R25214 vb.n83 vb.n82 54.344
R25215 vb.n100 vb.n99 54.344
R25216 vb.n190 vb.n189 51.092
R25217 vb.n180 vb.n178 50.947
R25218 vb.n72 vb.n71 47.551
R25219 vb.n111 vb.n110 47.551
R25220 vb.n178 vb.n4 46.314
R25221 vb.n177 vb.n176 44.423
R25222 vb.n16 vb.n15 44.155
R25223 vb.n165 vb.n164 44.155
R25224 vb.n61 vb.n60 40.758
R25225 vb.n122 vb.n121 40.758
R25226 vb.n27 vb.n26 37.362
R25227 vb.n154 vb.n153 37.362
R25228 vb.n50 vb.n49 33.965
R25229 vb.n133 vb.n132 33.965
R25230 vb.n38 vb.n37 30.568
R25231 vb.n143 vb.n142 30.568
R25232 vb.n39 vb.n38 27.172
R25233 vb.n144 vb.n143 27.172
R25234 vb.n193 vb.n192 24.1
R25235 vb.n49 vb.n48 23.775
R25236 vb.n132 vb.n131 23.775
R25237 vb.n28 vb.n27 20.379
R25238 vb.n155 vb.n154 20.379
R25239 vb.n60 vb.n59 16.982
R25240 vb.n121 vb.n120 16.982
R25241 vb.n17 vb.n16 13.586
R25242 vb.n166 vb.n165 13.586
R25243 vb.n91 vb.n90 13.176
R25244 vb.n71 vb.n70 10.189
R25245 vb.n110 vb.n109 10.189
R25246 vb.n172 vb.n171 9.3
R25247 vb.n161 vb.n160 9.3
R25248 vb.n150 vb.n149 9.3
R25249 vb.n139 vb.n138 9.3
R25250 vb.n128 vb.n127 9.3
R25251 vb.n117 vb.n116 9.3
R25252 vb.n106 vb.n105 9.3
R25253 vb.n94 vb.n93 9.3
R25254 vb.n87 vb.n86 9.3
R25255 vb.n76 vb.n75 9.3
R25256 vb.n65 vb.n64 9.3
R25257 vb.n54 vb.n53 9.3
R25258 vb.n43 vb.n42 9.3
R25259 vb.n32 vb.n31 9.3
R25260 vb.n21 vb.n20 9.3
R25261 vb.n10 vb.n9 9.3
R25262 vb.n8 vb.n7 9.3
R25263 vb.n12 vb.n11 9.3
R25264 vb.n19 vb.n18 9.3
R25265 vb.n18 vb.n17 9.3
R25266 vb.n23 vb.n22 9.3
R25267 vb.n30 vb.n29 9.3
R25268 vb.n29 vb.n28 9.3
R25269 vb.n34 vb.n33 9.3
R25270 vb.n41 vb.n40 9.3
R25271 vb.n40 vb.n39 9.3
R25272 vb.n45 vb.n44 9.3
R25273 vb.n52 vb.n51 9.3
R25274 vb.n51 vb.n50 9.3
R25275 vb.n56 vb.n55 9.3
R25276 vb.n63 vb.n62 9.3
R25277 vb.n62 vb.n61 9.3
R25278 vb.n67 vb.n66 9.3
R25279 vb.n74 vb.n73 9.3
R25280 vb.n73 vb.n72 9.3
R25281 vb.n78 vb.n77 9.3
R25282 vb.n85 vb.n84 9.3
R25283 vb.n84 vb.n83 9.3
R25284 vb.n89 vb.n88 9.3
R25285 vb.n92 vb.n91 9.3
R25286 vb.n102 vb.n101 9.3
R25287 vb.n101 vb.n100 9.3
R25288 vb.n104 vb.n103 9.3
R25289 vb.n113 vb.n112 9.3
R25290 vb.n112 vb.n111 9.3
R25291 vb.n115 vb.n114 9.3
R25292 vb.n124 vb.n123 9.3
R25293 vb.n123 vb.n122 9.3
R25294 vb.n126 vb.n125 9.3
R25295 vb.n135 vb.n134 9.3
R25296 vb.n134 vb.n133 9.3
R25297 vb.n137 vb.n136 9.3
R25298 vb.n146 vb.n145 9.3
R25299 vb.n145 vb.n144 9.3
R25300 vb.n148 vb.n147 9.3
R25301 vb.n157 vb.n156 9.3
R25302 vb.n156 vb.n155 9.3
R25303 vb.n159 vb.n158 9.3
R25304 vb.n168 vb.n167 9.3
R25305 vb.n167 vb.n166 9.3
R25306 vb.n170 vb.n169 9.3
R25307 vb.n175 vb.n174 9.3
R25308 vb.n4 vb 7.754
R25309 vb.n84 vb.n80 6.023
R25310 vb.n101 vb.n96 6.023
R25311 vb.n73 vb.n69 5.27
R25312 vb.n112 vb.n108 5.27
R25313 vb.n14 vb.n13 4.894
R25314 vb.n163 vb.n162 4.894
R25315 vb.n176 vb.n175 4.84
R25316 vb.n62 vb.n58 4.517
R25317 vb.n123 vb.n119 4.517
R25318 vb.n25 vb.n24 4.141
R25319 vb.n152 vb.n151 4.141
R25320 vb.n51 vb.n47 3.764
R25321 vb.n134 vb.n130 3.764
R25322 vb.n82 vb.n81 3.396
R25323 vb.n99 vb.n98 3.396
R25324 vb.n36 vb.n35 3.388
R25325 vb.n141 vb.n140 3.388
R25326 vb.n40 vb.n36 3.011
R25327 vb.n145 vb.n141 3.011
R25328 vb.n47 vb.n46 2.635
R25329 vb.n130 vb.n129 2.635
R25330 vb.n29 vb.n25 2.258
R25331 vb.n156 vb.n152 2.258
R25332 vb.n58 vb.n57 1.882
R25333 vb.n119 vb.n118 1.882
R25334 vb.n18 vb.n14 1.505
R25335 vb.n167 vb.n163 1.505
R25336 vb.n69 vb.n68 1.129
R25337 vb.n108 vb.n107 1.129
R25338 vb.n177 vb 0.853
R25339 vb.n7 vb.n6 0.851
R25340 vb.n174 vb.n173 0.851
R25341 vb.n80 vb.n79 0.376
R25342 vb.n96 vb.n95 0.376
R25343 vb.n8 vb.n5 0.19
R25344 vb.n92 vb.n89 0.19
R25345 vb.n19 vb.n12 0.144
R25346 vb.n30 vb.n23 0.144
R25347 vb.n41 vb.n34 0.144
R25348 vb.n52 vb.n45 0.144
R25349 vb.n63 vb.n56 0.144
R25350 vb.n74 vb.n67 0.144
R25351 vb.n85 vb.n78 0.144
R25352 vb.n104 vb.n102 0.144
R25353 vb.n115 vb.n113 0.144
R25354 vb.n126 vb.n124 0.144
R25355 vb.n137 vb.n135 0.144
R25356 vb.n148 vb.n146 0.144
R25357 vb.n159 vb.n157 0.144
R25358 vb.n170 vb.n168 0.144
R25359 vb.n87 vb.n85 0.043
R25360 vb.n102 vb.n94 0.043
R25361 vb.n12 vb.n10 0.04
R25362 vb.n172 vb.n170 0.04
R25363 vb.n76 vb.n74 0.038
R25364 vb.n113 vb.n106 0.038
R25365 vb.n23 vb.n21 0.035
R25366 vb.n161 vb.n159 0.035
R25367 vb.n65 vb.n63 0.032
R25368 vb.n124 vb.n117 0.032
R25369 vb.n34 vb.n32 0.029
R25370 vb.n150 vb.n148 0.029
R25371 vb.n54 vb.n52 0.027
R25372 vb.n135 vb.n128 0.027
R25373 vb.n45 vb.n43 0.024
R25374 vb.n139 vb.n137 0.024
R25375 vb.n43 vb.n41 0.021
R25376 vb.n146 vb.n139 0.021
R25377 vb.n56 vb.n54 0.019
R25378 vb.n128 vb.n126 0.019
R25379 vb.n32 vb.n30 0.016
R25380 vb.n157 vb.n150 0.016
R25381 vb.n67 vb.n65 0.013
R25382 vb.n117 vb.n115 0.013
R25383 vb.n21 vb.n19 0.01
R25384 vb.n168 vb.n161 0.01
R25385 vb.n78 vb.n76 0.008
R25386 vb.n106 vb.n104 0.008
R25387 vb.n10 vb.n8 0.005
R25388 vb.n175 vb.n172 0.005
R25389 vb.n89 vb.n87 0.002
R25390 vb.n94 vb.n92 0.002
R25391 va.n13 va 5667.83
R25392 va.n195 va.n194 791.384
R25393 va.n195 va 360.532
R25394 va.n249 va.t7 244.947
R25395 va.n14 va.n13 239.836
R25396 va.n243 va.t1 218.92
R25397 va.n2 va.t6 218.92
R25398 va.n240 va.t8 218.92
R25399 va.n1 va.t3 218.92
R25400 va.n237 va.t5 218.92
R25401 va.n0 va.t2 218.92
R25402 va.n234 va.t4 218.92
R25403 va.n230 va.t0 218.919
R25404 va.n109 va.n108 176.62
R25405 va.n235 va.n234 105.076
R25406 va.n233 va.n231 87.99
R25407 va.n250 va.n248 85.333
R25408 va.n248 va.n247 85.333
R25409 va.n247 va.n246 85.333
R25410 va.n246 va.n245 85.333
R25411 va.n245 va.n242 85.333
R25412 va.n242 va.n239 85.333
R25413 va.n239 va.n236 85.333
R25414 va.n236 va.n233 85.333
R25415 va.n238 va.n237 78.084
R25416 va.n250 va.n249 76
R25417 va.n248 va.n0 76
R25418 va.n247 va.n1 76
R25419 va.n246 va.n2 76
R25420 va.n245 va.n244 76
R25421 va.n242 va.n241 76
R25422 va.n239 va.n238 76
R25423 va.n236 va.n235 76
R25424 va.n233 va.n232 76
R25425 va.n12 va 73.93
R25426 va va.n250 68.266
R25427 va.n13 va.n12 58.619
R25428 va.n109 va.n107 54.344
R25429 va.n92 va.n91 54.344
R25430 va.n241 va.n240 51.092
R25431 va.n185 va.n184 50.948
R25432 va.n120 va.n119 47.551
R25433 va.n81 va.n80 47.551
R25434 va.n174 va.n173 44.155
R25435 va.n25 va.n24 44.155
R25436 va.n221 va.n220 41.786
R25437 va.n131 va.n130 40.758
R25438 va.n70 va.n69 40.758
R25439 va.n163 va.n162 37.362
R25440 va.n36 va.n35 37.362
R25441 va.n142 va.n141 33.965
R25442 va.n59 va.n58 33.965
R25443 va.n152 va.n151 30.568
R25444 va.n47 va.n46 30.568
R25445 va.n196 va.n195 29.778
R25446 va.n153 va.n152 27.172
R25447 va.n48 va.n47 27.172
R25448 va.n4 va.n3 24.204
R25449 va.n244 va.n243 24.1
R25450 va.n141 va.n140 23.775
R25451 va.n58 va.n57 23.775
R25452 va.n204 va.n201 21.438
R25453 va.n164 va.n163 20.379
R25454 va.n37 va.n36 20.379
R25455 va.n130 va.n129 16.982
R25456 va.n69 va.n68 16.982
R25457 va.n231 va.n230 16.194
R25458 va.n10 va 13.994
R25459 va.n175 va.n174 13.586
R25460 va.n26 va.n25 13.586
R25461 va.n100 va.n99 13.176
R25462 va.n231 va.n229 12.078
R25463 va.n119 va.n118 10.189
R25464 va.n80 va.n79 10.189
R25465 va.n19 va.n18 9.3
R25466 va.n30 va.n29 9.3
R25467 va.n41 va.n40 9.3
R25468 va.n52 va.n51 9.3
R25469 va.n63 va.n62 9.3
R25470 va.n74 va.n73 9.3
R25471 va.n85 va.n84 9.3
R25472 va.n96 va.n95 9.3
R25473 va.n103 va.n102 9.3
R25474 va.n115 va.n114 9.3
R25475 va.n126 va.n125 9.3
R25476 va.n137 va.n136 9.3
R25477 va.n148 va.n147 9.3
R25478 va.n159 va.n158 9.3
R25479 va.n170 va.n169 9.3
R25480 va.n188 va.n187 9.3
R25481 va.n187 va.n186 9.3
R25482 va.n17 va.n16 9.3
R25483 va.n21 va.n20 9.3
R25484 va.n28 va.n27 9.3
R25485 va.n27 va.n26 9.3
R25486 va.n32 va.n31 9.3
R25487 va.n39 va.n38 9.3
R25488 va.n38 va.n37 9.3
R25489 va.n43 va.n42 9.3
R25490 va.n50 va.n49 9.3
R25491 va.n49 va.n48 9.3
R25492 va.n54 va.n53 9.3
R25493 va.n61 va.n60 9.3
R25494 va.n60 va.n59 9.3
R25495 va.n65 va.n64 9.3
R25496 va.n72 va.n71 9.3
R25497 va.n71 va.n70 9.3
R25498 va.n76 va.n75 9.3
R25499 va.n83 va.n82 9.3
R25500 va.n82 va.n81 9.3
R25501 va.n87 va.n86 9.3
R25502 va.n94 va.n93 9.3
R25503 va.n93 va.n92 9.3
R25504 va.n98 va.n97 9.3
R25505 va.n101 va.n100 9.3
R25506 va.n111 va.n110 9.3
R25507 va.n110 va.n109 9.3
R25508 va.n113 va.n112 9.3
R25509 va.n122 va.n121 9.3
R25510 va.n121 va.n120 9.3
R25511 va.n124 va.n123 9.3
R25512 va.n133 va.n132 9.3
R25513 va.n132 va.n131 9.3
R25514 va.n135 va.n134 9.3
R25515 va.n144 va.n143 9.3
R25516 va.n143 va.n142 9.3
R25517 va.n146 va.n145 9.3
R25518 va.n155 va.n154 9.3
R25519 va.n154 va.n153 9.3
R25520 va.n157 va.n156 9.3
R25521 va.n166 va.n165 9.3
R25522 va.n165 va.n164 9.3
R25523 va.n168 va.n167 9.3
R25524 va.n177 va.n176 9.3
R25525 va.n176 va.n175 9.3
R25526 va.n179 va.n178 9.3
R25527 va.n181 va.n180 9.3
R25528 va.n197 va.n196 8.706
R25529 va.n186 va.n185 6.793
R25530 va.n110 va.n105 6.023
R25531 va.n93 va.n89 6.023
R25532 va.n183 va.n182 5.647
R25533 va.n193 va.n192 5.338
R25534 va.n121 va.n117 5.27
R25535 va.n82 va.n78 5.27
R25536 va.n172 va.n171 4.894
R25537 va.n23 va.n22 4.894
R25538 va.n17 va.n14 4.84
R25539 va.n204 va.n203 4.635
R25540 va.n12 va 4.547
R25541 va.n132 va.n128 4.517
R25542 va.n71 va.n67 4.517
R25543 va.n192 va.n191 4.374
R25544 va.n161 va.n160 4.141
R25545 va.n34 va.n33 4.141
R25546 va.n143 va.n139 3.764
R25547 va.n60 va.n56 3.764
R25548 va.n107 va.n106 3.396
R25549 va.n91 va.n90 3.396
R25550 va.n150 va.n149 3.388
R25551 va.n45 va.n44 3.388
R25552 va.n213 va.n212 3.186
R25553 va.n154 va.n150 3.011
R25554 va.n49 va.n45 3.011
R25555 va.n191 va.n190 2.635
R25556 va.n139 va.n138 2.635
R25557 va.n56 va.n55 2.635
R25558 va.n214 va.n213 2.325
R25559 va.n205 va.n204 2.325
R25560 va.n165 va.n161 2.258
R25561 va.n38 va.n34 2.258
R25562 va.n11 va.n10 2.116
R25563 va.n194 va 1.91
R25564 va.n128 va.n127 1.882
R25565 va.n67 va.n66 1.882
R25566 va.n194 va.n193 1.775
R25567 va.n212 va.n211 1.738
R25568 va.n193 va 1.676
R25569 va.n176 va.n172 1.505
R25570 va.n27 va.n23 1.505
R25571 va.n117 va.n116 1.129
R25572 va.n78 va.n77 1.129
R25573 va.n10 va 0.996
R25574 va.n11 va 0.995
R25575 va.n223 va.n221 0.885
R25576 va.n16 va.n15 0.851
R25577 va.n198 va.n9 0.775
R25578 va.n227 va.n226 0.775
R25579 va.n224 va.n223 0.775
R25580 va.n216 va.n215 0.775
R25581 va.n223 va.n222 0.774
R25582 va.n187 va.n183 0.752
R25583 va.n226 va.n225 0.7
R25584 va.n208 va 0.645
R25585 va.n219 va.n6 0.578
R25586 va.n228 va.n5 0.573
R25587 va.n105 va.n104 0.376
R25588 va.n89 va.n88 0.376
R25589 va va.n207 0.331
R25590 va.n205 va.n6 0.3
R25591 va.n206 va.n205 0.295
R25592 va.n203 va.n202 0.289
R25593 va.n5 va.n4 0.275
R25594 va.n215 va.n214 0.202
R25595 va.n214 va.n210 0.202
R25596 va.n9 va.n7 0.202
R25597 va.n101 va.n98 0.19
R25598 va.n189 va.n188 0.171
R25599 va.n179 va.n177 0.144
R25600 va.n168 va.n166 0.144
R25601 va.n157 va.n155 0.144
R25602 va.n146 va.n144 0.144
R25603 va.n135 va.n133 0.144
R25604 va.n124 va.n122 0.144
R25605 va.n113 va.n111 0.144
R25606 va.n94 va.n87 0.144
R25607 va.n83 va.n76 0.144
R25608 va.n72 va.n65 0.144
R25609 va.n61 va.n54 0.144
R25610 va.n50 va.n43 0.144
R25611 va.n39 va.n32 0.144
R25612 va.n28 va.n21 0.144
R25613 va.n215 va.n208 0.11
R25614 va.n210 va.n209 0.11
R25615 va.n9 va.n8 0.11
R25616 va.n196 va.n11 0.1
R25617 va.n111 va.n103 0.043
R25618 va.n96 va.n94 0.043
R25619 va.n181 va.n179 0.04
R25620 va.n21 va.n19 0.04
R25621 va.n122 va.n115 0.038
R25622 va.n85 va.n83 0.038
R25623 va.n170 va.n168 0.035
R25624 va.n32 va.n30 0.035
R25625 va.n133 va.n126 0.032
R25626 va.n74 va.n72 0.032
R25627 va.n159 va.n157 0.029
R25628 va.n43 va.n41 0.029
R25629 va.n144 va.n137 0.027
R25630 va.n63 va.n61 0.027
R25631 va.n192 va.n189 0.025
R25632 va.n148 va.n146 0.024
R25633 va.n54 va.n52 0.024
R25634 va.n155 va.n148 0.021
R25635 va.n52 va.n50 0.021
R25636 va.n227 va.n224 0.02
R25637 va.n224 va.n219 0.02
R25638 va.n137 va.n135 0.019
R25639 va.n65 va.n63 0.019
R25640 va.n228 va.n227 0.019
R25641 va.n207 va.n206 0.018
R25642 va.n166 va.n159 0.016
R25643 va.n41 va.n39 0.016
R25644 va.n218 va.n217 0.015
R25645 va.n200 va.n199 0.015
R25646 va.n126 va.n124 0.013
R25647 va.n76 va.n74 0.013
R25648 va.n177 va.n170 0.01
R25649 va.n30 va.n28 0.01
R25650 va.n115 va.n113 0.008
R25651 va.n87 va.n85 0.008
R25652 va.n188 va.n181 0.005
R25653 va.n19 va.n17 0.005
R25654 va.n219 va.n218 0.003
R25655 va.n103 va.n101 0.002
R25656 va.n98 va.n96 0.002
R25657 va.n229 va.n228 0.002
R25658 va.n216 va.n200 0.002
R25659 va.n199 va.n198 0.002
R25660 va.n217 va.n216 0.001
R25661 va.n198 va.n197 0.001
R25662 porst.n0 porst.t7 244.947
R25663 porst.n8 porst.t1 218.92
R25664 porst.n13 porst.t8 218.92
R25665 porst.n6 porst.t6 218.92
R25666 porst.n16 porst.t5 218.92
R25667 porst.n4 porst.t3 218.92
R25668 porst.n19 porst.t4 218.92
R25669 porst.n2 porst.t2 218.92
R25670 porst.n22 porst.t0 218.919
R25671 porst porst.n23 158.05
R25672 porst.n3 porst.n1 85.333
R25673 porst.n5 porst.n3 85.333
R25674 porst.n7 porst.n5 85.333
R25675 porst.n10 porst.n7 85.333
R25676 porst.n12 porst.n10 85.333
R25677 porst.n15 porst.n12 85.333
R25678 porst.n18 porst.n15 85.333
R25679 porst.n21 porst.n18 85.333
R25680 porst.n23 porst.n21 85.333
R25681 porst.n14 porst.n13 83.868
R25682 porst.n23 porst.n22 78.892
R25683 porst.n1 porst.n0 76
R25684 porst.n3 porst.n2 76
R25685 porst.n5 porst.n4 76
R25686 porst.n7 porst.n6 76
R25687 porst.n10 porst.n9 76
R25688 porst.n12 porst.n11 76
R25689 porst.n15 porst.n14 76
R25690 porst.n18 porst.n17 76
R25691 porst.n21 porst.n20 76
R25692 porst.n1 porst 68.266
R25693 porst.n17 porst.n16 56.876
R25694 porst.n20 porst.n19 29.884
R25695 porst.n9 porst.n8 24.1
R25696 sky130_asc_pfet_01v8_lvt_6_1/GATE.n81 sky130_asc_pfet_01v8_lvt_6_1/GATE.n80 875.047
R25697 sky130_asc_pfet_01v8_lvt_6_1/GATE.n203 sky130_asc_pfet_01v8_lvt_6_1/GATE.n202 239.836
R25698 sky130_asc_pfet_01v8_lvt_6_1/GATE.n74 sky130_asc_pfet_01v8_lvt_6_1/GATE.t12 222.22
R25699 sky130_asc_pfet_01v8_lvt_6_1/GATE.n34 sky130_asc_pfet_01v8_lvt_6_1/GATE.t10 222.22
R25700 sky130_asc_pfet_01v8_lvt_6_1/GATE.n205 sky130_asc_pfet_01v8_lvt_6_1/GATE.n204 195.413
R25701 sky130_asc_pfet_01v8_lvt_6_1/GATE.n204 sky130_asc_pfet_01v8_lvt_6_1/GATE.n203 195.413
R25702 sky130_asc_pfet_01v8_lvt_6_1/GATE.n66 sky130_asc_pfet_01v8_lvt_6_1/GATE.t16 166.1
R25703 sky130_asc_pfet_01v8_lvt_6_1/GATE.n26 sky130_asc_pfet_01v8_lvt_6_1/GATE.t2 166.1
R25704 sky130_asc_pfet_01v8_lvt_6_1/GATE.n71 sky130_asc_pfet_01v8_lvt_6_1/GATE.t17 166.1
R25705 sky130_asc_pfet_01v8_lvt_6_1/GATE.n60 sky130_asc_pfet_01v8_lvt_6_1/GATE.t15 166.1
R25706 sky130_asc_pfet_01v8_lvt_6_1/GATE.n24 sky130_asc_pfet_01v8_lvt_6_1/GATE.t4 166.1
R25707 sky130_asc_pfet_01v8_lvt_6_1/GATE.n31 sky130_asc_pfet_01v8_lvt_6_1/GATE.t0 166.1
R25708 sky130_asc_pfet_01v8_lvt_6_1/GATE.n69 sky130_asc_pfet_01v8_lvt_6_1/GATE.t13 166.1
R25709 sky130_asc_pfet_01v8_lvt_6_1/GATE.n35 sky130_asc_pfet_01v8_lvt_6_1/GATE.t8 166.1
R25710 sky130_asc_pfet_01v8_lvt_6_1/GATE.n75 sky130_asc_pfet_01v8_lvt_6_1/GATE.t14 166.1
R25711 sky130_asc_pfet_01v8_lvt_6_1/GATE.n36 sky130_asc_pfet_01v8_lvt_6_1/GATE.t6 166.1
R25712 sky130_asc_pfet_01v8_lvt_6_1/GATE.n67 sky130_asc_pfet_01v8_lvt_6_1/GATE.n66 126.284
R25713 sky130_asc_pfet_01v8_lvt_6_1/GATE.n77 sky130_asc_pfet_01v8_lvt_6_1/GATE.n74 122.204
R25714 sky130_asc_pfet_01v8_lvt_6_1/GATE.n38 sky130_asc_pfet_01v8_lvt_6_1/GATE.n34 122.204
R25715 sky130_asc_pfet_01v8_lvt_6_1/GATE.n71 sky130_asc_pfet_01v8_lvt_6_1/GATE.n70 100.256
R25716 sky130_asc_pfet_01v8_lvt_6_1/GATE.n32 sky130_asc_pfet_01v8_lvt_6_1/GATE.n31 100.256
R25717 sky130_asc_pfet_01v8_lvt_6_1/GATE.n81 sky130_asc_pfet_01v8_lvt_6_1/GATE 91.306
R25718 sky130_asc_pfet_01v8_lvt_6_1/GATE.n76 sky130_asc_pfet_01v8_lvt_6_1/GATE.n75 88.688
R25719 sky130_asc_pfet_01v8_lvt_6_1/GATE.n37 sky130_asc_pfet_01v8_lvt_6_1/GATE.n36 88.688
R25720 sky130_asc_pfet_01v8_lvt_6_1/GATE.n62 sky130_asc_pfet_01v8_lvt_6_1/GATE.n61 85.333
R25721 sky130_asc_pfet_01v8_lvt_6_1/GATE.n78 sky130_asc_pfet_01v8_lvt_6_1/GATE.n77 85.333
R25722 sky130_asc_pfet_01v8_lvt_6_1/GATE.n28 sky130_asc_pfet_01v8_lvt_6_1/GATE.n25 85.333
R25723 sky130_asc_pfet_01v8_lvt_6_1/GATE.n30 sky130_asc_pfet_01v8_lvt_6_1/GATE.n28 85.333
R25724 sky130_asc_pfet_01v8_lvt_6_1/GATE.n33 sky130_asc_pfet_01v8_lvt_6_1/GATE.n30 85.333
R25725 sky130_asc_pfet_01v8_lvt_6_1/GATE.n63 sky130_asc_pfet_01v8_lvt_6_1/GATE.n62 84.906
R25726 sky130_asc_pfet_01v8_lvt_6_1/GATE.n79 sky130_asc_pfet_01v8_lvt_6_1/GATE.n78 78.506
R25727 sky130_asc_pfet_01v8_lvt_6_1/GATE.n83 sky130_asc_pfet_01v8_lvt_6_1/GATE.n81 78.235
R25728 sky130_asc_pfet_01v8_lvt_6_1/GATE.n77 sky130_asc_pfet_01v8_lvt_6_1/GATE.n76 76
R25729 sky130_asc_pfet_01v8_lvt_6_1/GATE.n61 sky130_asc_pfet_01v8_lvt_6_1/GATE.n60 76
R25730 sky130_asc_pfet_01v8_lvt_6_1/GATE.n28 sky130_asc_pfet_01v8_lvt_6_1/GATE.n27 76
R25731 sky130_asc_pfet_01v8_lvt_6_1/GATE.n30 sky130_asc_pfet_01v8_lvt_6_1/GATE.n29 76
R25732 sky130_asc_pfet_01v8_lvt_6_1/GATE.n33 sky130_asc_pfet_01v8_lvt_6_1/GATE.n32 76
R25733 sky130_asc_pfet_01v8_lvt_6_1/GATE.n38 sky130_asc_pfet_01v8_lvt_6_1/GATE.n37 76
R25734 sky130_asc_pfet_01v8_lvt_6_1/GATE.n25 sky130_asc_pfet_01v8_lvt_6_1/GATE.n24 76
R25735 sky130_asc_pfet_01v8_lvt_6_1/GATE.n37 sky130_asc_pfet_01v8_lvt_6_1/GATE.n35 73.264
R25736 sky130_asc_pfet_01v8_lvt_6_1/GATE.n39 sky130_asc_pfet_01v8_lvt_6_1/GATE.n33 65.706
R25737 sky130_asc_pfet_01v8_lvt_6_1/GATE.n70 sky130_asc_pfet_01v8_lvt_6_1/GATE.n69 61.696
R25738 sky130_asc_pfet_01v8_lvt_6_1/GATE.n205 sky130_asc_pfet_01v8_lvt_6_1/GATE.t5 52.312
R25739 sky130_asc_pfet_01v8_lvt_6_1/GATE.n204 sky130_asc_pfet_01v8_lvt_6_1/GATE.n23 47.884
R25740 sky130_asc_pfet_01v8_lvt_6_1/GATE.n203 sky130_asc_pfet_01v8_lvt_6_1/GATE.n41 46.86
R25741 sky130_asc_pfet_01v8_lvt_6_1/GATE.n61 sky130_asc_pfet_01v8_lvt_6_1/GATE 46.08
R25742 sky130_asc_pfet_01v8_lvt_6_1/GATE.n25 sky130_asc_pfet_01v8_lvt_6_1/GATE 46.08
R25743 sky130_asc_pfet_01v8_lvt_6_1/GATE.n122 sky130_asc_pfet_01v8_lvt_6_1/GATE.n121 31.034
R25744 sky130_asc_pfet_01v8_lvt_6_1/GATE.n113 sky130_asc_pfet_01v8_lvt_6_1/GATE.n112 31.034
R25745 sky130_asc_pfet_01v8_lvt_6_1/GATE.n72 sky130_asc_pfet_01v8_lvt_6_1/GATE.n71 27.474
R25746 sky130_asc_pfet_01v8_lvt_6_1/GATE.n130 sky130_asc_pfet_01v8_lvt_6_1/GATE.n129 26.896
R25747 sky130_asc_pfet_01v8_lvt_6_1/GATE.n105 sky130_asc_pfet_01v8_lvt_6_1/GATE.n104 26.896
R25748 sky130_asc_pfet_01v8_lvt_6_1/GATE.n138 sky130_asc_pfet_01v8_lvt_6_1/GATE.n137 22.758
R25749 sky130_asc_pfet_01v8_lvt_6_1/GATE.n97 sky130_asc_pfet_01v8_lvt_6_1/GATE.n96 22.758
R25750 sky130_asc_pfet_01v8_lvt_6_1/GATE.n152 sky130_asc_pfet_01v8_lvt_6_1/GATE.n151 20.972
R25751 sky130_asc_pfet_01v8_lvt_6_1/GATE.n39 sky130_asc_pfet_01v8_lvt_6_1/GATE.n38 19.626
R25752 sky130_asc_pfet_01v8_lvt_6_1/GATE.n146 sky130_asc_pfet_01v8_lvt_6_1/GATE.n145 18.62
R25753 sky130_asc_pfet_01v8_lvt_6_1/GATE.n89 sky130_asc_pfet_01v8_lvt_6_1/GATE.n88 18.62
R25754 sky130_asc_pfet_01v8_lvt_6_1/GATE.n147 sky130_asc_pfet_01v8_lvt_6_1/GATE.n146 16.551
R25755 sky130_asc_pfet_01v8_lvt_6_1/GATE.n90 sky130_asc_pfet_01v8_lvt_6_1/GATE.n89 16.551
R25756 sky130_asc_pfet_01v8_lvt_6_1/GATE.n173 sky130_asc_pfet_01v8_lvt_6_1/GATE.n172 13.176
R25757 sky130_asc_pfet_01v8_lvt_6_1/GATE.n139 sky130_asc_pfet_01v8_lvt_6_1/GATE.n138 12.413
R25758 sky130_asc_pfet_01v8_lvt_6_1/GATE.n98 sky130_asc_pfet_01v8_lvt_6_1/GATE.n97 12.413
R25759 sky130_asc_pfet_01v8_lvt_6_1/GATE.n73 sky130_asc_pfet_01v8_lvt_6_1/GATE.n72 9.3
R25760 sky130_asc_pfet_01v8_lvt_6_1/GATE.n22 sky130_asc_pfet_01v8_lvt_6_1/GATE.n149 9.3
R25761 sky130_asc_pfet_01v8_lvt_6_1/GATE.n18 sky130_asc_pfet_01v8_lvt_6_1/GATE.n141 9.3
R25762 sky130_asc_pfet_01v8_lvt_6_1/GATE.n12 sky130_asc_pfet_01v8_lvt_6_1/GATE.n133 9.3
R25763 sky130_asc_pfet_01v8_lvt_6_1/GATE.n8 sky130_asc_pfet_01v8_lvt_6_1/GATE.n125 9.3
R25764 sky130_asc_pfet_01v8_lvt_6_1/GATE.n7 sky130_asc_pfet_01v8_lvt_6_1/GATE.n109 9.3
R25765 sky130_asc_pfet_01v8_lvt_6_1/GATE.n11 sky130_asc_pfet_01v8_lvt_6_1/GATE.n101 9.3
R25766 sky130_asc_pfet_01v8_lvt_6_1/GATE.n17 sky130_asc_pfet_01v8_lvt_6_1/GATE.n93 9.3
R25767 sky130_asc_pfet_01v8_lvt_6_1/GATE.n21 sky130_asc_pfet_01v8_lvt_6_1/GATE.n85 9.3
R25768 sky130_asc_pfet_01v8_lvt_6_1/GATE.n21 sky130_asc_pfet_01v8_lvt_6_1/GATE.n84 9.3
R25769 sky130_asc_pfet_01v8_lvt_6_1/GATE.n21 sky130_asc_pfet_01v8_lvt_6_1/GATE.n91 9.3
R25770 sky130_asc_pfet_01v8_lvt_6_1/GATE.n91 sky130_asc_pfet_01v8_lvt_6_1/GATE.n90 9.3
R25771 sky130_asc_pfet_01v8_lvt_6_1/GATE.n17 sky130_asc_pfet_01v8_lvt_6_1/GATE.n92 9.3
R25772 sky130_asc_pfet_01v8_lvt_6_1/GATE.n17 sky130_asc_pfet_01v8_lvt_6_1/GATE.n99 9.3
R25773 sky130_asc_pfet_01v8_lvt_6_1/GATE.n99 sky130_asc_pfet_01v8_lvt_6_1/GATE.n98 9.3
R25774 sky130_asc_pfet_01v8_lvt_6_1/GATE.n11 sky130_asc_pfet_01v8_lvt_6_1/GATE.n100 9.3
R25775 sky130_asc_pfet_01v8_lvt_6_1/GATE.n11 sky130_asc_pfet_01v8_lvt_6_1/GATE.n107 9.3
R25776 sky130_asc_pfet_01v8_lvt_6_1/GATE.n107 sky130_asc_pfet_01v8_lvt_6_1/GATE.n106 9.3
R25777 sky130_asc_pfet_01v8_lvt_6_1/GATE.n7 sky130_asc_pfet_01v8_lvt_6_1/GATE.n108 9.3
R25778 sky130_asc_pfet_01v8_lvt_6_1/GATE.n7 sky130_asc_pfet_01v8_lvt_6_1/GATE.n115 9.3
R25779 sky130_asc_pfet_01v8_lvt_6_1/GATE.n115 sky130_asc_pfet_01v8_lvt_6_1/GATE.n114 9.3
R25780 sky130_asc_pfet_01v8_lvt_6_1/GATE.n8 sky130_asc_pfet_01v8_lvt_6_1/GATE.n124 9.3
R25781 sky130_asc_pfet_01v8_lvt_6_1/GATE.n124 sky130_asc_pfet_01v8_lvt_6_1/GATE.n123 9.3
R25782 sky130_asc_pfet_01v8_lvt_6_1/GATE.n8 sky130_asc_pfet_01v8_lvt_6_1/GATE.n126 9.3
R25783 sky130_asc_pfet_01v8_lvt_6_1/GATE.n12 sky130_asc_pfet_01v8_lvt_6_1/GATE.n132 9.3
R25784 sky130_asc_pfet_01v8_lvt_6_1/GATE.n132 sky130_asc_pfet_01v8_lvt_6_1/GATE.n131 9.3
R25785 sky130_asc_pfet_01v8_lvt_6_1/GATE.n12 sky130_asc_pfet_01v8_lvt_6_1/GATE.n134 9.3
R25786 sky130_asc_pfet_01v8_lvt_6_1/GATE.n18 sky130_asc_pfet_01v8_lvt_6_1/GATE.n140 9.3
R25787 sky130_asc_pfet_01v8_lvt_6_1/GATE.n140 sky130_asc_pfet_01v8_lvt_6_1/GATE.n139 9.3
R25788 sky130_asc_pfet_01v8_lvt_6_1/GATE.n18 sky130_asc_pfet_01v8_lvt_6_1/GATE.n142 9.3
R25789 sky130_asc_pfet_01v8_lvt_6_1/GATE.n22 sky130_asc_pfet_01v8_lvt_6_1/GATE.n148 9.3
R25790 sky130_asc_pfet_01v8_lvt_6_1/GATE.n148 sky130_asc_pfet_01v8_lvt_6_1/GATE.n147 9.3
R25791 sky130_asc_pfet_01v8_lvt_6_1/GATE.n22 sky130_asc_pfet_01v8_lvt_6_1/GATE.n150 9.3
R25792 sky130_asc_pfet_01v8_lvt_6_1/GATE.n10 sky130_asc_pfet_01v8_lvt_6_1/GATE.n154 9.3
R25793 sky130_asc_pfet_01v8_lvt_6_1/GATE.n16 sky130_asc_pfet_01v8_lvt_6_1/GATE.n156 9.3
R25794 sky130_asc_pfet_01v8_lvt_6_1/GATE.n20 sky130_asc_pfet_01v8_lvt_6_1/GATE.n158 9.3
R25795 sky130_asc_pfet_01v8_lvt_6_1/GATE.n3 sky130_asc_pfet_01v8_lvt_6_1/GATE.n160 9.3
R25796 sky130_asc_pfet_01v8_lvt_6_1/GATE.n14 sky130_asc_pfet_01v8_lvt_6_1/GATE.n163 9.3
R25797 sky130_asc_pfet_01v8_lvt_6_1/GATE.n1 sky130_asc_pfet_01v8_lvt_6_1/GATE.n166 9.3
R25798 sky130_asc_pfet_01v8_lvt_6_1/GATE.n6 sky130_asc_pfet_01v8_lvt_6_1/GATE.n170 9.3
R25799 sky130_asc_pfet_01v8_lvt_6_1/GATE.n5 sky130_asc_pfet_01v8_lvt_6_1/GATE.n174 9.3
R25800 sky130_asc_pfet_01v8_lvt_6_1/GATE.n0 sky130_asc_pfet_01v8_lvt_6_1/GATE.n178 9.3
R25801 sky130_asc_pfet_01v8_lvt_6_1/GATE.n13 sky130_asc_pfet_01v8_lvt_6_1/GATE.n182 9.3
R25802 sky130_asc_pfet_01v8_lvt_6_1/GATE.n2 sky130_asc_pfet_01v8_lvt_6_1/GATE.n186 9.3
R25803 sky130_asc_pfet_01v8_lvt_6_1/GATE.n19 sky130_asc_pfet_01v8_lvt_6_1/GATE.n190 9.3
R25804 sky130_asc_pfet_01v8_lvt_6_1/GATE.n15 sky130_asc_pfet_01v8_lvt_6_1/GATE.n194 9.3
R25805 sky130_asc_pfet_01v8_lvt_6_1/GATE.n9 sky130_asc_pfet_01v8_lvt_6_1/GATE.n198 9.3
R25806 sky130_asc_pfet_01v8_lvt_6_1/GATE.n4 sky130_asc_pfet_01v8_lvt_6_1/GATE.n201 9.3
R25807 sky130_asc_pfet_01v8_lvt_6_1/GATE.n9 sky130_asc_pfet_01v8_lvt_6_1/GATE.n197 9.3
R25808 sky130_asc_pfet_01v8_lvt_6_1/GATE.n15 sky130_asc_pfet_01v8_lvt_6_1/GATE.n193 9.3
R25809 sky130_asc_pfet_01v8_lvt_6_1/GATE.n19 sky130_asc_pfet_01v8_lvt_6_1/GATE.n189 9.3
R25810 sky130_asc_pfet_01v8_lvt_6_1/GATE.n2 sky130_asc_pfet_01v8_lvt_6_1/GATE.n185 9.3
R25811 sky130_asc_pfet_01v8_lvt_6_1/GATE.n13 sky130_asc_pfet_01v8_lvt_6_1/GATE.n181 9.3
R25812 sky130_asc_pfet_01v8_lvt_6_1/GATE.n0 sky130_asc_pfet_01v8_lvt_6_1/GATE.n177 9.3
R25813 sky130_asc_pfet_01v8_lvt_6_1/GATE.n5 sky130_asc_pfet_01v8_lvt_6_1/GATE.n173 9.3
R25814 sky130_asc_pfet_01v8_lvt_6_1/GATE.n6 sky130_asc_pfet_01v8_lvt_6_1/GATE.n171 9.3
R25815 sky130_asc_pfet_01v8_lvt_6_1/GATE.n1 sky130_asc_pfet_01v8_lvt_6_1/GATE.n167 9.3
R25816 sky130_asc_pfet_01v8_lvt_6_1/GATE.n14 sky130_asc_pfet_01v8_lvt_6_1/GATE.n164 9.3
R25817 sky130_asc_pfet_01v8_lvt_6_1/GATE.n3 sky130_asc_pfet_01v8_lvt_6_1/GATE.n161 9.3
R25818 sky130_asc_pfet_01v8_lvt_6_1/GATE.n20 sky130_asc_pfet_01v8_lvt_6_1/GATE.n159 9.3
R25819 sky130_asc_pfet_01v8_lvt_6_1/GATE.n16 sky130_asc_pfet_01v8_lvt_6_1/GATE.n157 9.3
R25820 sky130_asc_pfet_01v8_lvt_6_1/GATE.n10 sky130_asc_pfet_01v8_lvt_6_1/GATE.n155 9.3
R25821 sky130_asc_pfet_01v8_lvt_6_1/GATE.n152 sky130_asc_pfet_01v8_lvt_6_1/GATE.n153 9.3
R25822 sky130_asc_pfet_01v8_lvt_6_1/GATE.n9 sky130_asc_pfet_01v8_lvt_6_1/GATE.n200 9.3
R25823 sky130_asc_pfet_01v8_lvt_6_1/GATE.n15 sky130_asc_pfet_01v8_lvt_6_1/GATE.n196 9.3
R25824 sky130_asc_pfet_01v8_lvt_6_1/GATE.n19 sky130_asc_pfet_01v8_lvt_6_1/GATE.n192 9.3
R25825 sky130_asc_pfet_01v8_lvt_6_1/GATE.n2 sky130_asc_pfet_01v8_lvt_6_1/GATE.n188 9.3
R25826 sky130_asc_pfet_01v8_lvt_6_1/GATE.n13 sky130_asc_pfet_01v8_lvt_6_1/GATE.n184 9.3
R25827 sky130_asc_pfet_01v8_lvt_6_1/GATE.n0 sky130_asc_pfet_01v8_lvt_6_1/GATE.n180 9.3
R25828 sky130_asc_pfet_01v8_lvt_6_1/GATE.n5 sky130_asc_pfet_01v8_lvt_6_1/GATE.n176 9.3
R25829 sky130_asc_pfet_01v8_lvt_6_1/GATE.n6 sky130_asc_pfet_01v8_lvt_6_1/GATE.n169 9.3
R25830 sky130_asc_pfet_01v8_lvt_6_1/GATE.n1 sky130_asc_pfet_01v8_lvt_6_1/GATE.n165 9.3
R25831 sky130_asc_pfet_01v8_lvt_6_1/GATE.n14 sky130_asc_pfet_01v8_lvt_6_1/GATE.n162 9.3
R25832 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n43 8.896
R25833 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n51 8.885
R25834 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n45 8.875
R25835 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n49 8.864
R25836 sky130_asc_pfet_01v8_lvt_6_1/GATE.n117 sky130_asc_pfet_01v8_lvt_6_1/GATE.n116 8.855
R25837 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n46 8.853
R25838 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n47 8.843
R25839 sky130_asc_pfet_01v8_lvt_6_1/GATE.n131 sky130_asc_pfet_01v8_lvt_6_1/GATE.n130 8.275
R25840 sky130_asc_pfet_01v8_lvt_6_1/GATE.n106 sky130_asc_pfet_01v8_lvt_6_1/GATE.n105 8.275
R25841 sky130_asc_pfet_01v8_lvt_6_1/GATE.n66 sky130_asc_pfet_01v8_lvt_6_1/GATE.n65 7.712
R25842 sky130_asc_pfet_01v8_lvt_6_1/GATE.n27 sky130_asc_pfet_01v8_lvt_6_1/GATE.n26 7.712
R25843 sky130_asc_pfet_01v8_lvt_6_1/GATE.n72 sky130_asc_pfet_01v8_lvt_6_1/GATE.n68 7.23
R25844 sky130_asc_pfet_01v8_lvt_6_1/GATE.n41 sky130_asc_pfet_01v8_lvt_6_1/GATE.n39 6.553
R25845 sky130_asc_pfet_01v8_lvt_6_1/GATE.n151 sky130_asc_pfet_01v8_lvt_6_1/GATE.n59 6.084
R25846 sky130_asc_pfet_01v8_lvt_6_1/GATE.n120 sky130_asc_pfet_01v8_lvt_6_1/GATE.n119 5.647
R25847 sky130_asc_pfet_01v8_lvt_6_1/GATE.n111 sky130_asc_pfet_01v8_lvt_6_1/GATE.n110 5.647
R25848 sky130_asc_pfet_01v8_lvt_6_1/GATE.n202 sky130_asc_pfet_01v8_lvt_6_1/GATE.n58 5.417
R25849 sky130_asc_pfet_01v8_lvt_6_1/GATE.n58 sky130_asc_pfet_01v8_lvt_6_1/GATE.n57 5.382
R25850 sky130_asc_pfet_01v8_lvt_6_1/GATE.n54 sky130_asc_pfet_01v8_lvt_6_1/GATE.n53 5.379
R25851 sky130_asc_pfet_01v8_lvt_6_1/GATE.n128 sky130_asc_pfet_01v8_lvt_6_1/GATE.n127 4.894
R25852 sky130_asc_pfet_01v8_lvt_6_1/GATE.n103 sky130_asc_pfet_01v8_lvt_6_1/GATE.n102 4.894
R25853 sky130_asc_pfet_01v8_lvt_6_1/GATE.n202 sky130_asc_pfet_01v8_lvt_6_1/GATE.n4 4.84
R25854 sky130_asc_pfet_01v8_lvt_6_1/GATE.n118 sky130_asc_pfet_01v8_lvt_6_1/GATE.n117 4.65
R25855 sky130_asc_pfet_01v8_lvt_6_1/GATE.n23 sky130_asc_pfet_01v8_lvt_6_1/GATE.t3 4.428
R25856 sky130_asc_pfet_01v8_lvt_6_1/GATE.n23 sky130_asc_pfet_01v8_lvt_6_1/GATE.t1 4.428
R25857 sky130_asc_pfet_01v8_lvt_6_1/GATE.n40 sky130_asc_pfet_01v8_lvt_6_1/GATE.t9 4.428
R25858 sky130_asc_pfet_01v8_lvt_6_1/GATE.n40 sky130_asc_pfet_01v8_lvt_6_1/GATE.t7 4.428
R25859 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.t11 4.428
R25860 sky130_asc_pfet_01v8_lvt_6_1/GATE.n136 sky130_asc_pfet_01v8_lvt_6_1/GATE.n135 4.141
R25861 sky130_asc_pfet_01v8_lvt_6_1/GATE.n95 sky130_asc_pfet_01v8_lvt_6_1/GATE.n94 4.141
R25862 sky130_asc_pfet_01v8_lvt_6_1/GATE.n123 sky130_asc_pfet_01v8_lvt_6_1/GATE.n122 4.137
R25863 sky130_asc_pfet_01v8_lvt_6_1/GATE.n114 sky130_asc_pfet_01v8_lvt_6_1/GATE.n113 4.137
R25864 sky130_asc_pfet_01v8_lvt_6_1/GATE.n83 sky130_asc_pfet_01v8_lvt_6_1/GATE.n82 3.954
R25865 sky130_asc_pfet_01v8_lvt_6_1/GATE.n144 sky130_asc_pfet_01v8_lvt_6_1/GATE.n143 3.388
R25866 sky130_asc_pfet_01v8_lvt_6_1/GATE.n87 sky130_asc_pfet_01v8_lvt_6_1/GATE.n86 3.388
R25867 sky130_asc_pfet_01v8_lvt_6_1/GATE.n73 sky130_asc_pfet_01v8_lvt_6_1/GATE.n64 3.2
R25868 sky130_asc_pfet_01v8_lvt_6_1/GATE.n80 sky130_asc_pfet_01v8_lvt_6_1/GATE.n73 3.2
R25869 sky130_asc_pfet_01v8_lvt_6_1/GATE.n148 sky130_asc_pfet_01v8_lvt_6_1/GATE.n144 3.011
R25870 sky130_asc_pfet_01v8_lvt_6_1/GATE.n91 sky130_asc_pfet_01v8_lvt_6_1/GATE.n87 3.011
R25871 sky130_asc_pfet_01v8_lvt_6_1/GATE.n140 sky130_asc_pfet_01v8_lvt_6_1/GATE.n136 2.258
R25872 sky130_asc_pfet_01v8_lvt_6_1/GATE.n99 sky130_asc_pfet_01v8_lvt_6_1/GATE.n95 2.258
R25873 sky130_asc_pfet_01v8_lvt_6_1/GATE.n21 sky130_asc_pfet_01v8_lvt_6_1/GATE.n83 2.249
R25874 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 sky130_asc_pfet_01v8_lvt_6_1/GATE.n54 1.844
R25875 sky130_asc_pfet_01v8_lvt_6_1/GATE.n58 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 1.844
R25876 sky130_asc_pfet_01v8_lvt_6_1/GATE.n132 sky130_asc_pfet_01v8_lvt_6_1/GATE.n128 1.505
R25877 sky130_asc_pfet_01v8_lvt_6_1/GATE.n107 sky130_asc_pfet_01v8_lvt_6_1/GATE.n103 1.505
R25878 sky130_asc_pfet_01v8_lvt_6_1/GATE.n41 sky130_asc_pfet_01v8_lvt_6_1/GATE.n40 1.023
R25879 sky130_asc_pfet_01v8_lvt_6_1/GATE.n68 sky130_asc_pfet_01v8_lvt_6_1/GATE.n67 0.964
R25880 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_pfet_01v8_lvt_6_1/GATE.n205 0.853
R25881 sky130_asc_pfet_01v8_lvt_6_1/GATE.n124 sky130_asc_pfet_01v8_lvt_6_1/GATE.n120 0.752
R25882 sky130_asc_pfet_01v8_lvt_6_1/GATE.n115 sky130_asc_pfet_01v8_lvt_6_1/GATE.n111 0.752
R25883 sky130_asc_pfet_01v8_lvt_6_1/GATE.n53 sky130_asc_pfet_01v8_lvt_6_1/GATE.n52 0.752
R25884 sky130_asc_pfet_01v8_lvt_6_1/GATE.n57 sky130_asc_pfet_01v8_lvt_6_1/GATE.n56 0.752
R25885 sky130_asc_pfet_01v8_lvt_6_1/GATE.n64 sky130_asc_pfet_01v8_lvt_6_1/GATE.n63 0.426
R25886 sky130_asc_pfet_01v8_lvt_6_1/GATE.n80 sky130_asc_pfet_01v8_lvt_6_1/GATE.n79 0.426
R25887 sky130_asc_pfet_01v8_lvt_6_1/GATE.n6 sky130_asc_pfet_01v8_lvt_6_1/GATE.n1 0.235
R25888 sky130_asc_pfet_01v8_lvt_6_1/GATE.n12 sky130_asc_pfet_01v8_lvt_6_1/GATE.n8 0.234
R25889 sky130_asc_pfet_01v8_lvt_6_1/GATE.n7 sky130_asc_pfet_01v8_lvt_6_1/GATE.n11 0.234
R25890 sky130_asc_pfet_01v8_lvt_6_1/GATE.n4 sky130_asc_pfet_01v8_lvt_6_1/GATE.n9 0.234
R25891 sky130_asc_pfet_01v8_lvt_6_1/GATE.n8 sky130_asc_pfet_01v8_lvt_6_1/GATE.n118 0.19
R25892 sky130_asc_pfet_01v8_lvt_6_1/GATE.n118 sky130_asc_pfet_01v8_lvt_6_1/GATE.n7 0.19
R25893 sky130_asc_pfet_01v8_lvt_6_1/GATE.n5 sky130_asc_pfet_01v8_lvt_6_1/GATE.n6 0.19
R25894 sky130_asc_pfet_01v8_lvt_6_1/GATE.n14 sky130_asc_pfet_01v8_lvt_6_1/GATE.n3 0.19
R25895 sky130_asc_pfet_01v8_lvt_6_1/GATE.n19 sky130_asc_pfet_01v8_lvt_6_1/GATE.n2 0.19
R25896 sky130_asc_pfet_01v8_lvt_6_1/GATE.n13 sky130_asc_pfet_01v8_lvt_6_1/GATE.n0 0.19
R25897 sky130_asc_pfet_01v8_lvt_6_1/GATE.n22 sky130_asc_pfet_01v8_lvt_6_1/GATE.n18 0.189
R25898 sky130_asc_pfet_01v8_lvt_6_1/GATE.n17 sky130_asc_pfet_01v8_lvt_6_1/GATE.n21 0.189
R25899 sky130_asc_pfet_01v8_lvt_6_1/GATE.n3 sky130_asc_pfet_01v8_lvt_6_1/GATE.n20 0.189
R25900 sky130_asc_pfet_01v8_lvt_6_1/GATE.n15 sky130_asc_pfet_01v8_lvt_6_1/GATE.n19 0.189
R25901 sky130_asc_pfet_01v8_lvt_6_1/GATE.n18 sky130_asc_pfet_01v8_lvt_6_1/GATE.n12 0.189
R25902 sky130_asc_pfet_01v8_lvt_6_1/GATE.n11 sky130_asc_pfet_01v8_lvt_6_1/GATE.n17 0.189
R25903 sky130_asc_pfet_01v8_lvt_6_1/GATE.n20 sky130_asc_pfet_01v8_lvt_6_1/GATE.n16 0.189
R25904 sky130_asc_pfet_01v8_lvt_6_1/GATE.n9 sky130_asc_pfet_01v8_lvt_6_1/GATE.n15 0.189
R25905 sky130_asc_pfet_01v8_lvt_6_1/GATE.n1 sky130_asc_pfet_01v8_lvt_6_1/GATE.n14 0.189
R25906 sky130_asc_pfet_01v8_lvt_6_1/GATE.n2 sky130_asc_pfet_01v8_lvt_6_1/GATE.n13 0.189
R25907 sky130_asc_pfet_01v8_lvt_6_1/GATE.n16 sky130_asc_pfet_01v8_lvt_6_1/GATE.n10 0.189
R25908 sky130_asc_pfet_01v8_lvt_6_1/GATE.n0 sky130_asc_pfet_01v8_lvt_6_1/GATE.n5 0.189
R25909 sky130_asc_pfet_01v8_lvt_6_1/GATE.n176 sky130_asc_pfet_01v8_lvt_6_1/GATE.n175 0.189
R25910 sky130_asc_pfet_01v8_lvt_6_1/GATE.n169 sky130_asc_pfet_01v8_lvt_6_1/GATE.n168 0.188
R25911 sky130_asc_pfet_01v8_lvt_6_1/GATE.n180 sky130_asc_pfet_01v8_lvt_6_1/GATE.n179 0.178
R25912 sky130_asc_pfet_01v8_lvt_6_1/GATE.n184 sky130_asc_pfet_01v8_lvt_6_1/GATE.n183 0.166
R25913 sky130_asc_pfet_01v8_lvt_6_1/GATE.n151 sky130_asc_pfet_01v8_lvt_6_1/GATE.n22 0.163
R25914 sky130_asc_pfet_01v8_lvt_6_1/GATE.n188 sky130_asc_pfet_01v8_lvt_6_1/GATE.n187 0.155
R25915 sky130_asc_pfet_01v8_lvt_6_1/GATE.n49 sky130_asc_pfet_01v8_lvt_6_1/GATE.n48 0.155
R25916 sky130_asc_pfet_01v8_lvt_6_1/GATE.n192 sky130_asc_pfet_01v8_lvt_6_1/GATE.n191 0.144
R25917 sky130_asc_pfet_01v8_lvt_6_1/GATE.n10 sky130_asc_pfet_01v8_lvt_6_1/GATE.n152 0.144
R25918 sky130_asc_pfet_01v8_lvt_6_1/GATE.n45 sky130_asc_pfet_01v8_lvt_6_1/GATE.n44 0.144
R25919 sky130_asc_pfet_01v8_lvt_6_1/GATE.n196 sky130_asc_pfet_01v8_lvt_6_1/GATE.n195 0.133
R25920 sky130_asc_pfet_01v8_lvt_6_1/GATE.n51 sky130_asc_pfet_01v8_lvt_6_1/GATE.n50 0.132
R25921 sky130_asc_pfet_01v8_lvt_6_1/GATE.n200 sky130_asc_pfet_01v8_lvt_6_1/GATE.n199 0.121
R25922 sky130_asc_pfet_01v8_lvt_6_1/GATE.n43 sky130_asc_pfet_01v8_lvt_6_1/GATE.n42 0.121
C0 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.68fF
C1 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin 1.25fF
C2 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# VDD 0.00fF
C3 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.28fF
C4 sky130_asc_res_xhigh_po_2p85_1_17/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin -0.31fF
C5 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.29fF
C6 sky130_asc_res_xhigh_po_2p85_1_1/Rin vbg 0.03fF
C7 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.54fF
C8 sky130_asc_res_xhigh_po_2p85_1_9/Rin VDD 3.19fF
C9 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.20fF
C10 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.12fF
C11 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.69fF
C12 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.33fF
C13 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.45fF
C14 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.03fF
C15 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.45fF
C16 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# vb 1.19fF
C17 sky130_asc_res_xhigh_po_2p85_1_17/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.03fF
C18 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.15fF
C19 va sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.67fF
C20 sky130_asc_res_xhigh_po_2p85_1_11/Rin vbg 0.03fF
C21 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.29fF
C22 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.03fF
C23 sky130_asc_res_xhigh_po_2p85_1_21/Rin VDD 0.32fF
C24 sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.20fF
C25 sky130_asc_res_xhigh_po_2p85_1_24/Rin va 1.28fF
C26 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_2_0/Rin 1.27fF
C27 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.04fF
C28 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.52fF
C29 sky130_asc_cap_mim_m3_1_4/Cout VDD 2.40fF
C30 porst VDD 0.74fF
C31 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb 0.45fF
C32 sky130_asc_nfet_01v8_lvt_1_1/GATE va 2.67fF
C33 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.64fF
C34 sky130_asc_res_xhigh_po_2p85_1_19/Rin VDD 0.21fF
C35 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.20fF
C36 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.76fF
C37 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.20fF
C38 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.06fF
C39 sky130_asc_res_xhigh_po_2p85_1_29/Rin VDD 0.85fF
C40 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.09fF
C41 sky130_asc_res_xhigh_po_2p85_1_6/Rin VDD 0.11fF
C42 sky130_asc_nfet_01v8_lvt_1_1/GATE vb 0.21fF
C43 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.48fF
C44 va sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.04fF
C45 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.11fF
C46 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.03fF
C47 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VDD 6.46fF
C48 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.56fF
C49 sky130_asc_res_xhigh_po_2p85_1_4/Rin VDD 0.12fF
C50 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.45fF
C51 sky130_asc_pfet_01v8_lvt_6_1/GATE vb 1.33fF
C52 sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.57fF
C53 sky130_asc_res_xhigh_po_2p85_1_23/Rin vb 0.04fF
C54 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.31fF
C55 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.53fF
C56 sky130_asc_res_xhigh_po_2p85_2_0/Rin VDD 0.89fF
C57 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.31fF
C58 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.20fF
C59 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.06fF
C60 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin 1.27fF
C61 sky130_asc_res_xhigh_po_2p85_1_9/Rin vb 0.03fF
C62 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# 0.59fF
C63 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.20fF
C64 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rin 3.42fF
C65 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.67fF
C66 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# 0.27fF
C67 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 1.20fF
C68 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.49fF
C69 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.15fF
C70 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.46fF
C71 sky130_asc_res_xhigh_po_2p85_1_13/Rin VDD 1.32fF
C72 sky130_asc_cap_mim_m3_1_4/Cout va 0.14fF
C73 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_2_0/Rin 1.92fF
C74 sky130_asc_res_xhigh_po_2p85_1_26/Rin VDD 4.52fF
C75 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.45fF
C76 sky130_asc_res_xhigh_po_2p85_1_7/Rin VDD 1.36fF
C77 sky130_asc_res_xhigh_po_2p85_1_19/Rout VDD 0.32fF
C78 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.10fF
C79 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.61fF
C80 sky130_asc_res_xhigh_po_2p85_1_5/Rin vbg 0.03fF
C81 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.08fF
C82 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.20fF
C83 sky130_asc_cap_mim_m3_1_4/Cout vb 1.46fF
C84 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.20fF
C85 vbg sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.03fF
C86 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.15fF
C87 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.20fF
C88 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.20fF
C89 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.03fF
C90 sky130_asc_res_xhigh_po_2p85_2_1/Rin VDD 0.11fF
C91 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.45fF
C92 sky130_asc_nfet_01v8_lvt_1_1/DRAIN va -0.09fF
C93 sky130_asc_res_xhigh_po_2p85_1_15/Rin VDD 8.78fF
C94 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.51fF
C95 va sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.04fF
C96 sky130_asc_res_xhigh_po_2p85_1_12/Rin VDD 0.80fF
C97 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.20fF
C98 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# 0.20fF
C99 sky130_asc_res_xhigh_po_2p85_1_18/Rin VDD 3.54fF
C100 va VDD 3.88fF
C101 sky130_asc_cap_mim_m3_1_4/Cout vbg 0.17fF
C102 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.20fF
C103 sky130_asc_res_xhigh_po_2p85_1_1/Rin VDD 2.00fF
C104 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_pfet_01v8_lvt_6_1/GATE 0.01fF
C105 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_res_xhigh_po_2p85_1_23/Rin 1.11fF
C106 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 6.50fF
C107 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.53fF
C108 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.03fF
C109 vb sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.04fF
C110 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.03fF
C111 va sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.03fF
C112 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_12/Rin 2.11fF
C113 vb VDD 5.18fF
C114 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.05fF
C115 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.29fF
C116 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.20fF
C117 sky130_asc_res_xhigh_po_2p85_1_11/Rin VDD 0.24fF
C118 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# sky130_asc_pfet_01v8_lvt_6_1/GATE 0.26fF
C119 vb sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.04fF
C120 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.03fF
C121 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.23fF
C122 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# va 0.23fF
C123 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.63fF
C124 sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.21fF
C125 sky130_asc_res_xhigh_po_2p85_1_19/Rout vb 0.51fF
C126 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_nfet_01v8_lvt_1_1/GATE 3.17fF
C127 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.03fF
C128 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.46fF
C129 sky130_asc_res_xhigh_po_2p85_1_15/Rin va 0.36fF
C130 vbg VDD 4.03fF
C131 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# vb 0.20fF
C132 sky130_asc_res_xhigh_po_2p85_1_10/Rin vb -0.29fF
C133 sky130_asc_res_xhigh_po_2p85_1_3/Rin vbg 0.03fF
C134 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.03fF
C135 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_pfet_01v8_lvt_6_1/GATE 0.27fF
C136 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# va 0.33fF
C137 sky130_asc_res_xhigh_po_2p85_1_15/Rin vb 0.45fF
C138 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_23/Rin 1.40fF
C139 sky130_asc_res_xhigh_po_2p85_1_25/Rin VDD 2.10fF
C140 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# vbg 0.20fF
C141 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.00fF
C142 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.46fF
C143 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.31fF
C144 sky130_asc_res_xhigh_po_2p85_1_14/Rin VDD 1.07fF
C145 vb sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.04fF
C146 sky130_asc_res_xhigh_po_2p85_1_17/Rin VDD 0.89fF
C147 sky130_asc_res_xhigh_po_2p85_1_27/Rin VDD 0.11fF
C148 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.33fF
C149 sky130_asc_res_xhigh_po_2p85_1_18/Rin vb 0.03fF
C150 va vb 0.04fF
C151 sky130_asc_res_xhigh_po_2p85_1_2/Rin VDD 0.11fF
C152 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.90fF
C153 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 1.35fF
C154 sky130_asc_res_xhigh_po_2p85_1_24/Rin VDD 1.11fF
C155 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.03fF
C156 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.45fF
C157 sky130_asc_nfet_01v8_lvt_1_1/GATE VDD 1.75fF
C158 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin 1.86fF
C159 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.36fF
C160 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/GATE 0.29fF
C161 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.03fF
C162 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.49fF
C163 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.31fF
C164 sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.20fF
C165 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.36fF
C166 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.29fF
C167 sky130_asc_res_xhigh_po_2p85_1_22/Rin VDD 0.11fF
C168 sky130_asc_cap_mim_m3_1_4/Cout porst 0.18fF
C169 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.22fF
C170 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.03fF
C171 sky130_asc_res_xhigh_po_2p85_1_5/Rin VDD 0.11fF
C172 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.16fF
C173 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD 3.23fF
C174 sky130_asc_res_xhigh_po_2p85_1_23/Rin VDD 2.69fF
C175 VDD VSS 1243.13fF
C176 porst VSS 35.60fF
C177 sky130_asc_res_xhigh_po_2p85_1_6/Rin VSS 2.95fF
C178 sky130_asc_res_xhigh_po_2p85_1_12/Rin VSS 5.85fF
C179 sky130_asc_res_xhigh_po_2p85_1_7/Rin VSS 6.02fF
C180 sky130_asc_res_xhigh_po_2p85_1_2/Rin VSS 2.74fF
C181 sky130_asc_res_xhigh_po_2p85_1_13/Rin VSS 2.53fF
C182 sky130_asc_res_xhigh_po_2p85_1_14/Rin VSS 3.52fF
C183 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS 9.87fF
C184 sky130_asc_res_xhigh_po_2p85_1_19/Rin VSS 3.51fF
C185 vb VSS 47.07fF
C186 sky130_asc_res_xhigh_po_2p85_1_18/Rin VSS 3.88fF
C187 sky130_asc_res_xhigh_po_2p85_1_9/Rin VSS 4.42fF
C188 sky130_asc_res_xhigh_po_2p85_1_10/Rin VSS 3.56fF
C189 sky130_asc_res_xhigh_po_2p85_1_22/Rin VSS 2.81fF
C190 sky130_asc_res_xhigh_po_2p85_1_23/Rin VSS 6.28fF
C191 sky130_asc_res_xhigh_po_2p85_1_28/Rin VSS 7.25fF
C192 sky130_asc_res_xhigh_po_2p85_1_26/Rin VSS 4.82fF
C193 sky130_asc_res_xhigh_po_2p85_1_27/Rin VSS 3.96fF
C194 sky130_asc_res_xhigh_po_2p85_1_21/Rin VSS 12.18fF
C195 vbg VSS 27.55fF
C196 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS 11.17fF
C197 sky130_asc_pfet_01v8_lvt_6_1/GATE.n0 VSS 0.01fF $ **FLOATING
C198 sky130_asc_pfet_01v8_lvt_6_1/GATE.n1 VSS 0.01fF $ **FLOATING
C199 sky130_asc_pfet_01v8_lvt_6_1/GATE.n2 VSS 0.01fF $ **FLOATING
C200 sky130_asc_pfet_01v8_lvt_6_1/GATE.n3 VSS 0.01fF $ **FLOATING
C201 sky130_asc_pfet_01v8_lvt_6_1/GATE.n4 VSS 0.02fF $ **FLOATING
C202 sky130_asc_pfet_01v8_lvt_6_1/GATE.n5 VSS 0.01fF $ **FLOATING
C203 sky130_asc_pfet_01v8_lvt_6_1/GATE.n6 VSS 0.01fF $ **FLOATING
C204 sky130_asc_pfet_01v8_lvt_6_1/GATE.n7 VSS 0.01fF $ **FLOATING
C205 sky130_asc_pfet_01v8_lvt_6_1/GATE.n8 VSS 0.01fF $ **FLOATING
C206 sky130_asc_pfet_01v8_lvt_6_1/GATE.n9 VSS 0.01fF $ **FLOATING
C207 sky130_asc_pfet_01v8_lvt_6_1/GATE.n10 VSS 0.01fF $ **FLOATING
C208 sky130_asc_pfet_01v8_lvt_6_1/GATE.n11 VSS 0.01fF $ **FLOATING
C209 sky130_asc_pfet_01v8_lvt_6_1/GATE.n12 VSS 0.01fF $ **FLOATING
C210 sky130_asc_pfet_01v8_lvt_6_1/GATE.n13 VSS 0.01fF $ **FLOATING
C211 sky130_asc_pfet_01v8_lvt_6_1/GATE.n14 VSS 0.01fF $ **FLOATING
C212 sky130_asc_pfet_01v8_lvt_6_1/GATE.n15 VSS 0.01fF $ **FLOATING
C213 sky130_asc_pfet_01v8_lvt_6_1/GATE.n16 VSS 0.01fF $ **FLOATING
C214 sky130_asc_pfet_01v8_lvt_6_1/GATE.n17 VSS 0.01fF $ **FLOATING
C215 sky130_asc_pfet_01v8_lvt_6_1/GATE.n18 VSS 0.01fF $ **FLOATING
C216 sky130_asc_pfet_01v8_lvt_6_1/GATE.n19 VSS 0.01fF $ **FLOATING
C217 sky130_asc_pfet_01v8_lvt_6_1/GATE.n20 VSS 0.01fF $ **FLOATING
C218 sky130_asc_pfet_01v8_lvt_6_1/GATE.n21 VSS 0.02fF $ **FLOATING
C219 sky130_asc_pfet_01v8_lvt_6_1/GATE.n22 VSS 0.01fF $ **FLOATING
C220 sky130_asc_pfet_01v8_lvt_6_1/GATE.t5 VSS 0.52fF
C221 sky130_asc_pfet_01v8_lvt_6_1/GATE.t3 VSS 0.06fF
C222 sky130_asc_pfet_01v8_lvt_6_1/GATE.t1 VSS 0.06fF
C223 sky130_asc_pfet_01v8_lvt_6_1/GATE.n23 VSS 0.45fF $ **FLOATING
C224 sky130_asc_pfet_01v8_lvt_6_1/GATE.t4 VSS 1.45fF
C225 sky130_asc_pfet_01v8_lvt_6_1/GATE.n24 VSS 0.26fF $ **FLOATING
C226 sky130_asc_pfet_01v8_lvt_6_1/GATE.n25 VSS 0.06fF $ **FLOATING
C227 sky130_asc_pfet_01v8_lvt_6_1/GATE.t2 VSS 1.45fF
C228 sky130_asc_pfet_01v8_lvt_6_1/GATE.n26 VSS 0.33fF $ **FLOATING
C229 sky130_asc_pfet_01v8_lvt_6_1/GATE.n27 VSS 0.05fF $ **FLOATING
C230 sky130_asc_pfet_01v8_lvt_6_1/GATE.n28 VSS 0.08fF $ **FLOATING
C231 sky130_asc_pfet_01v8_lvt_6_1/GATE.n29 VSS 0.05fF $ **FLOATING
C232 sky130_asc_pfet_01v8_lvt_6_1/GATE.n30 VSS 0.08fF $ **FLOATING
C233 sky130_asc_pfet_01v8_lvt_6_1/GATE.t0 VSS 1.45fF
C234 sky130_asc_pfet_01v8_lvt_6_1/GATE.n31 VSS 0.33fF $ **FLOATING
C235 sky130_asc_pfet_01v8_lvt_6_1/GATE.n32 VSS 0.05fF $ **FLOATING
C236 sky130_asc_pfet_01v8_lvt_6_1/GATE.n33 VSS 0.07fF $ **FLOATING
C237 sky130_asc_pfet_01v8_lvt_6_1/GATE.t10 VSS 1.56fF
C238 sky130_asc_pfet_01v8_lvt_6_1/GATE.n34 VSS 0.44fF $ **FLOATING
C239 sky130_asc_pfet_01v8_lvt_6_1/GATE.t8 VSS 1.45fF
C240 sky130_asc_pfet_01v8_lvt_6_1/GATE.n35 VSS 0.33fF $ **FLOATING
C241 sky130_asc_pfet_01v8_lvt_6_1/GATE.t6 VSS 1.45fF
C242 sky130_asc_pfet_01v8_lvt_6_1/GATE.n36 VSS 0.35fF $ **FLOATING
C243 sky130_asc_pfet_01v8_lvt_6_1/GATE.n37 VSS 0.05fF $ **FLOATING
C244 sky130_asc_pfet_01v8_lvt_6_1/GATE.n38 VSS 0.08fF $ **FLOATING
C245 sky130_asc_pfet_01v8_lvt_6_1/GATE.n39 VSS 0.06fF $ **FLOATING
C246 sky130_asc_pfet_01v8_lvt_6_1/GATE.t9 VSS 0.06fF
C247 sky130_asc_pfet_01v8_lvt_6_1/GATE.t7 VSS 0.06fF
C248 sky130_asc_pfet_01v8_lvt_6_1/GATE.n40 VSS 0.30fF $ **FLOATING
C249 sky130_asc_pfet_01v8_lvt_6_1/GATE.n41 VSS 0.16fF $ **FLOATING
C250 sky130_asc_pfet_01v8_lvt_6_1/GATE.t11 VSS 0.06fF
C251 sky130_asc_pfet_01v8_lvt_6_1/GATE.n42 VSS 0.00fF $ **FLOATING
C252 sky130_asc_pfet_01v8_lvt_6_1/GATE.n43 VSS 0.00fF $ **FLOATING
C253 sky130_asc_pfet_01v8_lvt_6_1/GATE.n44 VSS 0.00fF $ **FLOATING
C254 sky130_asc_pfet_01v8_lvt_6_1/GATE.n45 VSS 0.00fF $ **FLOATING
C255 sky130_asc_pfet_01v8_lvt_6_1/GATE.n46 VSS 0.00fF $ **FLOATING
C256 sky130_asc_pfet_01v8_lvt_6_1/GATE.n47 VSS 0.00fF $ **FLOATING
C257 sky130_asc_pfet_01v8_lvt_6_1/GATE.n48 VSS 0.00fF $ **FLOATING
C258 sky130_asc_pfet_01v8_lvt_6_1/GATE.n49 VSS 0.00fF $ **FLOATING
C259 sky130_asc_pfet_01v8_lvt_6_1/GATE.n50 VSS 0.00fF $ **FLOATING
C260 sky130_asc_pfet_01v8_lvt_6_1/GATE.n51 VSS 0.00fF $ **FLOATING
C261 sky130_asc_pfet_01v8_lvt_6_1/GATE.n52 VSS 0.00fF $ **FLOATING
C262 sky130_asc_pfet_01v8_lvt_6_1/GATE.n53 VSS 0.00fF $ **FLOATING
C263 sky130_asc_pfet_01v8_lvt_6_1/GATE.n54 VSS 0.00fF $ **FLOATING
C264 sky130_asc_pfet_01v8_lvt_6_1/GATE.n55 VSS 0.18fF $ **FLOATING
C265 sky130_asc_pfet_01v8_lvt_6_1/GATE.n56 VSS 0.00fF $ **FLOATING
C266 sky130_asc_pfet_01v8_lvt_6_1/GATE.n57 VSS 0.00fF $ **FLOATING
C267 sky130_asc_pfet_01v8_lvt_6_1/GATE.n58 VSS 0.00fF $ **FLOATING
C268 sky130_asc_pfet_01v8_lvt_6_1/GATE.n59 VSS 0.02fF $ **FLOATING
C269 sky130_asc_pfet_01v8_lvt_6_1/GATE.t15 VSS 1.45fF
C270 sky130_asc_pfet_01v8_lvt_6_1/GATE.n60 VSS 0.26fF $ **FLOATING
C271 sky130_asc_pfet_01v8_lvt_6_1/GATE.n61 VSS 0.06fF $ **FLOATING
C272 sky130_asc_pfet_01v8_lvt_6_1/GATE.n62 VSS 0.08fF $ **FLOATING
C273 sky130_asc_pfet_01v8_lvt_6_1/GATE.n63 VSS 0.04fF $ **FLOATING
C274 sky130_asc_pfet_01v8_lvt_6_1/GATE.n64 VSS 0.00fF $ **FLOATING
C275 sky130_asc_pfet_01v8_lvt_6_1/GATE.n65 VSS 0.05fF $ **FLOATING
C276 sky130_asc_pfet_01v8_lvt_6_1/GATE.t16 VSS 1.45fF
C277 sky130_asc_pfet_01v8_lvt_6_1/GATE.n66 VSS 0.33fF $ **FLOATING
C278 sky130_asc_pfet_01v8_lvt_6_1/GATE.n67 VSS 0.04fF $ **FLOATING
C279 sky130_asc_pfet_01v8_lvt_6_1/GATE.n68 VSS 0.00fF $ **FLOATING
C280 sky130_asc_pfet_01v8_lvt_6_1/GATE.t13 VSS 1.45fF
C281 sky130_asc_pfet_01v8_lvt_6_1/GATE.n69 VSS 0.33fF $ **FLOATING
C282 sky130_asc_pfet_01v8_lvt_6_1/GATE.n70 VSS 0.05fF $ **FLOATING
C283 sky130_asc_pfet_01v8_lvt_6_1/GATE.t17 VSS 1.45fF
C284 sky130_asc_pfet_01v8_lvt_6_1/GATE.n71 VSS 0.33fF $ **FLOATING
C285 sky130_asc_pfet_01v8_lvt_6_1/GATE.n72 VSS 0.01fF $ **FLOATING
C286 sky130_asc_pfet_01v8_lvt_6_1/GATE.n73 VSS 0.00fF $ **FLOATING
C287 sky130_asc_pfet_01v8_lvt_6_1/GATE.t12 VSS 1.56fF
C288 sky130_asc_pfet_01v8_lvt_6_1/GATE.n74 VSS 0.44fF $ **FLOATING
C289 sky130_asc_pfet_01v8_lvt_6_1/GATE.t14 VSS 1.45fF
C290 sky130_asc_pfet_01v8_lvt_6_1/GATE.n75 VSS 0.35fF $ **FLOATING
C291 sky130_asc_pfet_01v8_lvt_6_1/GATE.n76 VSS 0.05fF $ **FLOATING
C292 sky130_asc_pfet_01v8_lvt_6_1/GATE.n77 VSS 0.11fF $ **FLOATING
C293 sky130_asc_pfet_01v8_lvt_6_1/GATE.n78 VSS 0.07fF $ **FLOATING
C294 sky130_asc_pfet_01v8_lvt_6_1/GATE.n79 VSS 0.04fF $ **FLOATING
C295 sky130_asc_pfet_01v8_lvt_6_1/GATE.n80 VSS 1.36fF $ **FLOATING
C296 sky130_asc_pfet_01v8_lvt_6_1/GATE.n81 VSS 1.06fF $ **FLOATING
C297 sky130_asc_pfet_01v8_lvt_6_1/GATE.n82 VSS 0.02fF $ **FLOATING
C298 sky130_asc_pfet_01v8_lvt_6_1/GATE.n83 VSS 0.02fF $ **FLOATING
C299 sky130_asc_pfet_01v8_lvt_6_1/GATE.n84 VSS 0.00fF $ **FLOATING
C300 sky130_asc_pfet_01v8_lvt_6_1/GATE.n85 VSS 0.00fF $ **FLOATING
C301 sky130_asc_pfet_01v8_lvt_6_1/GATE.n86 VSS 0.00fF $ **FLOATING
C302 sky130_asc_pfet_01v8_lvt_6_1/GATE.n87 VSS 0.00fF $ **FLOATING
C303 sky130_asc_pfet_01v8_lvt_6_1/GATE.n88 VSS 0.01fF $ **FLOATING
C304 sky130_asc_pfet_01v8_lvt_6_1/GATE.n89 VSS 0.00fF $ **FLOATING
C305 sky130_asc_pfet_01v8_lvt_6_1/GATE.n90 VSS 0.01fF $ **FLOATING
C306 sky130_asc_pfet_01v8_lvt_6_1/GATE.n91 VSS 0.00fF $ **FLOATING
C307 sky130_asc_pfet_01v8_lvt_6_1/GATE.n92 VSS 0.00fF $ **FLOATING
C308 sky130_asc_pfet_01v8_lvt_6_1/GATE.n93 VSS 0.00fF $ **FLOATING
C309 sky130_asc_pfet_01v8_lvt_6_1/GATE.n94 VSS 0.00fF $ **FLOATING
C310 sky130_asc_pfet_01v8_lvt_6_1/GATE.n95 VSS 0.00fF $ **FLOATING
C311 sky130_asc_pfet_01v8_lvt_6_1/GATE.n96 VSS 0.01fF $ **FLOATING
C312 sky130_asc_pfet_01v8_lvt_6_1/GATE.n97 VSS 0.00fF $ **FLOATING
C313 sky130_asc_pfet_01v8_lvt_6_1/GATE.n98 VSS 0.01fF $ **FLOATING
C314 sky130_asc_pfet_01v8_lvt_6_1/GATE.n99 VSS 0.00fF $ **FLOATING
C315 sky130_asc_pfet_01v8_lvt_6_1/GATE.n100 VSS 0.00fF $ **FLOATING
C316 sky130_asc_pfet_01v8_lvt_6_1/GATE.n101 VSS 0.00fF $ **FLOATING
C317 sky130_asc_pfet_01v8_lvt_6_1/GATE.n102 VSS 0.00fF $ **FLOATING
C318 sky130_asc_pfet_01v8_lvt_6_1/GATE.n103 VSS 0.00fF $ **FLOATING
C319 sky130_asc_pfet_01v8_lvt_6_1/GATE.n104 VSS 0.01fF $ **FLOATING
C320 sky130_asc_pfet_01v8_lvt_6_1/GATE.n105 VSS 0.00fF $ **FLOATING
C321 sky130_asc_pfet_01v8_lvt_6_1/GATE.n106 VSS 0.01fF $ **FLOATING
C322 sky130_asc_pfet_01v8_lvt_6_1/GATE.n107 VSS 0.00fF $ **FLOATING
C323 sky130_asc_pfet_01v8_lvt_6_1/GATE.n108 VSS 0.00fF $ **FLOATING
C324 sky130_asc_pfet_01v8_lvt_6_1/GATE.n109 VSS 0.00fF $ **FLOATING
C325 sky130_asc_pfet_01v8_lvt_6_1/GATE.n110 VSS 0.00fF $ **FLOATING
C326 sky130_asc_pfet_01v8_lvt_6_1/GATE.n111 VSS 0.00fF $ **FLOATING
C327 sky130_asc_pfet_01v8_lvt_6_1/GATE.n112 VSS 0.01fF $ **FLOATING
C328 sky130_asc_pfet_01v8_lvt_6_1/GATE.n113 VSS 0.00fF $ **FLOATING
C329 sky130_asc_pfet_01v8_lvt_6_1/GATE.n114 VSS 0.01fF $ **FLOATING
C330 sky130_asc_pfet_01v8_lvt_6_1/GATE.n115 VSS 0.00fF $ **FLOATING
C331 sky130_asc_pfet_01v8_lvt_6_1/GATE.n116 VSS 0.01fF $ **FLOATING
C332 sky130_asc_pfet_01v8_lvt_6_1/GATE.n117 VSS 0.01fF $ **FLOATING
C333 sky130_asc_pfet_01v8_lvt_6_1/GATE.n118 VSS 0.01fF $ **FLOATING
C334 sky130_asc_pfet_01v8_lvt_6_1/GATE.n119 VSS 0.00fF $ **FLOATING
C335 sky130_asc_pfet_01v8_lvt_6_1/GATE.n120 VSS 0.00fF $ **FLOATING
C336 sky130_asc_pfet_01v8_lvt_6_1/GATE.n121 VSS 0.01fF $ **FLOATING
C337 sky130_asc_pfet_01v8_lvt_6_1/GATE.n122 VSS 0.00fF $ **FLOATING
C338 sky130_asc_pfet_01v8_lvt_6_1/GATE.n123 VSS 0.01fF $ **FLOATING
C339 sky130_asc_pfet_01v8_lvt_6_1/GATE.n124 VSS 0.00fF $ **FLOATING
C340 sky130_asc_pfet_01v8_lvt_6_1/GATE.n125 VSS 0.00fF $ **FLOATING
C341 sky130_asc_pfet_01v8_lvt_6_1/GATE.n126 VSS 0.00fF $ **FLOATING
C342 sky130_asc_pfet_01v8_lvt_6_1/GATE.n127 VSS 0.00fF $ **FLOATING
C343 sky130_asc_pfet_01v8_lvt_6_1/GATE.n128 VSS 0.00fF $ **FLOATING
C344 sky130_asc_pfet_01v8_lvt_6_1/GATE.n129 VSS 0.01fF $ **FLOATING
C345 sky130_asc_pfet_01v8_lvt_6_1/GATE.n130 VSS 0.00fF $ **FLOATING
C346 sky130_asc_pfet_01v8_lvt_6_1/GATE.n131 VSS 0.01fF $ **FLOATING
C347 sky130_asc_pfet_01v8_lvt_6_1/GATE.n132 VSS 0.00fF $ **FLOATING
C348 sky130_asc_pfet_01v8_lvt_6_1/GATE.n133 VSS 0.00fF $ **FLOATING
C349 sky130_asc_pfet_01v8_lvt_6_1/GATE.n134 VSS 0.00fF $ **FLOATING
C350 sky130_asc_pfet_01v8_lvt_6_1/GATE.n135 VSS 0.00fF $ **FLOATING
C351 sky130_asc_pfet_01v8_lvt_6_1/GATE.n136 VSS 0.00fF $ **FLOATING
C352 sky130_asc_pfet_01v8_lvt_6_1/GATE.n137 VSS 0.01fF $ **FLOATING
C353 sky130_asc_pfet_01v8_lvt_6_1/GATE.n138 VSS 0.00fF $ **FLOATING
C354 sky130_asc_pfet_01v8_lvt_6_1/GATE.n139 VSS 0.01fF $ **FLOATING
C355 sky130_asc_pfet_01v8_lvt_6_1/GATE.n140 VSS 0.00fF $ **FLOATING
C356 sky130_asc_pfet_01v8_lvt_6_1/GATE.n141 VSS 0.00fF $ **FLOATING
C357 sky130_asc_pfet_01v8_lvt_6_1/GATE.n142 VSS 0.00fF $ **FLOATING
C358 sky130_asc_pfet_01v8_lvt_6_1/GATE.n143 VSS 0.00fF $ **FLOATING
C359 sky130_asc_pfet_01v8_lvt_6_1/GATE.n144 VSS 0.00fF $ **FLOATING
C360 sky130_asc_pfet_01v8_lvt_6_1/GATE.n145 VSS 0.01fF $ **FLOATING
C361 sky130_asc_pfet_01v8_lvt_6_1/GATE.n146 VSS 0.00fF $ **FLOATING
C362 sky130_asc_pfet_01v8_lvt_6_1/GATE.n147 VSS 0.01fF $ **FLOATING
C363 sky130_asc_pfet_01v8_lvt_6_1/GATE.n148 VSS 0.00fF $ **FLOATING
C364 sky130_asc_pfet_01v8_lvt_6_1/GATE.n149 VSS 0.00fF $ **FLOATING
C365 sky130_asc_pfet_01v8_lvt_6_1/GATE.n150 VSS 0.00fF $ **FLOATING
C366 sky130_asc_pfet_01v8_lvt_6_1/GATE.n151 VSS 0.23fF $ **FLOATING
C367 sky130_asc_pfet_01v8_lvt_6_1/GATE.n152 VSS 0.23fF $ **FLOATING
C368 sky130_asc_pfet_01v8_lvt_6_1/GATE.n153 VSS 0.00fF $ **FLOATING
C369 sky130_asc_pfet_01v8_lvt_6_1/GATE.n154 VSS 0.00fF $ **FLOATING
C370 sky130_asc_pfet_01v8_lvt_6_1/GATE.n155 VSS 0.00fF $ **FLOATING
C371 sky130_asc_pfet_01v8_lvt_6_1/GATE.n156 VSS 0.00fF $ **FLOATING
C372 sky130_asc_pfet_01v8_lvt_6_1/GATE.n157 VSS 0.00fF $ **FLOATING
C373 sky130_asc_pfet_01v8_lvt_6_1/GATE.n158 VSS 0.00fF $ **FLOATING
C374 sky130_asc_pfet_01v8_lvt_6_1/GATE.n159 VSS 0.00fF $ **FLOATING
C375 sky130_asc_pfet_01v8_lvt_6_1/GATE.n160 VSS 0.00fF $ **FLOATING
C376 sky130_asc_pfet_01v8_lvt_6_1/GATE.n161 VSS 0.00fF $ **FLOATING
C377 sky130_asc_pfet_01v8_lvt_6_1/GATE.n162 VSS 0.00fF $ **FLOATING
C378 sky130_asc_pfet_01v8_lvt_6_1/GATE.n163 VSS 0.00fF $ **FLOATING
C379 sky130_asc_pfet_01v8_lvt_6_1/GATE.n164 VSS 0.00fF $ **FLOATING
C380 sky130_asc_pfet_01v8_lvt_6_1/GATE.n165 VSS 0.00fF $ **FLOATING
C381 sky130_asc_pfet_01v8_lvt_6_1/GATE.n166 VSS 0.00fF $ **FLOATING
C382 sky130_asc_pfet_01v8_lvt_6_1/GATE.n167 VSS 0.00fF $ **FLOATING
C383 sky130_asc_pfet_01v8_lvt_6_1/GATE.n168 VSS 0.00fF $ **FLOATING
C384 sky130_asc_pfet_01v8_lvt_6_1/GATE.n169 VSS 0.00fF $ **FLOATING
C385 sky130_asc_pfet_01v8_lvt_6_1/GATE.n170 VSS 0.00fF $ **FLOATING
C386 sky130_asc_pfet_01v8_lvt_6_1/GATE.n171 VSS 0.00fF $ **FLOATING
C387 sky130_asc_pfet_01v8_lvt_6_1/GATE.n172 VSS 0.00fF $ **FLOATING
C388 sky130_asc_pfet_01v8_lvt_6_1/GATE.n173 VSS 0.00fF $ **FLOATING
C389 sky130_asc_pfet_01v8_lvt_6_1/GATE.n174 VSS 0.00fF $ **FLOATING
C390 sky130_asc_pfet_01v8_lvt_6_1/GATE.n175 VSS 0.00fF $ **FLOATING
C391 sky130_asc_pfet_01v8_lvt_6_1/GATE.n176 VSS 0.00fF $ **FLOATING
C392 sky130_asc_pfet_01v8_lvt_6_1/GATE.n177 VSS 0.00fF $ **FLOATING
C393 sky130_asc_pfet_01v8_lvt_6_1/GATE.n178 VSS 0.00fF $ **FLOATING
C394 sky130_asc_pfet_01v8_lvt_6_1/GATE.n179 VSS 0.00fF $ **FLOATING
C395 sky130_asc_pfet_01v8_lvt_6_1/GATE.n180 VSS 0.00fF $ **FLOATING
C396 sky130_asc_pfet_01v8_lvt_6_1/GATE.n181 VSS 0.00fF $ **FLOATING
C397 sky130_asc_pfet_01v8_lvt_6_1/GATE.n182 VSS 0.00fF $ **FLOATING
C398 sky130_asc_pfet_01v8_lvt_6_1/GATE.n183 VSS 0.00fF $ **FLOATING
C399 sky130_asc_pfet_01v8_lvt_6_1/GATE.n184 VSS 0.00fF $ **FLOATING
C400 sky130_asc_pfet_01v8_lvt_6_1/GATE.n185 VSS 0.00fF $ **FLOATING
C401 sky130_asc_pfet_01v8_lvt_6_1/GATE.n186 VSS 0.00fF $ **FLOATING
C402 sky130_asc_pfet_01v8_lvt_6_1/GATE.n187 VSS 0.00fF $ **FLOATING
C403 sky130_asc_pfet_01v8_lvt_6_1/GATE.n188 VSS 0.00fF $ **FLOATING
C404 sky130_asc_pfet_01v8_lvt_6_1/GATE.n189 VSS 0.00fF $ **FLOATING
C405 sky130_asc_pfet_01v8_lvt_6_1/GATE.n190 VSS 0.00fF $ **FLOATING
C406 sky130_asc_pfet_01v8_lvt_6_1/GATE.n191 VSS 0.00fF $ **FLOATING
C407 sky130_asc_pfet_01v8_lvt_6_1/GATE.n192 VSS 0.00fF $ **FLOATING
C408 sky130_asc_pfet_01v8_lvt_6_1/GATE.n193 VSS 0.00fF $ **FLOATING
C409 sky130_asc_pfet_01v8_lvt_6_1/GATE.n194 VSS 0.00fF $ **FLOATING
C410 sky130_asc_pfet_01v8_lvt_6_1/GATE.n195 VSS 0.00fF $ **FLOATING
C411 sky130_asc_pfet_01v8_lvt_6_1/GATE.n196 VSS 0.00fF $ **FLOATING
C412 sky130_asc_pfet_01v8_lvt_6_1/GATE.n197 VSS 0.00fF $ **FLOATING
C413 sky130_asc_pfet_01v8_lvt_6_1/GATE.n198 VSS 0.00fF $ **FLOATING
C414 sky130_asc_pfet_01v8_lvt_6_1/GATE.n199 VSS 0.00fF $ **FLOATING
C415 sky130_asc_pfet_01v8_lvt_6_1/GATE.n200 VSS 0.00fF $ **FLOATING
C416 sky130_asc_pfet_01v8_lvt_6_1/GATE.n201 VSS 0.00fF $ **FLOATING
C417 sky130_asc_pfet_01v8_lvt_6_1/GATE.n202 VSS 0.10fF $ **FLOATING
C418 sky130_asc_pfet_01v8_lvt_6_1/GATE.n203 VSS 0.20fF $ **FLOATING
C419 sky130_asc_pfet_01v8_lvt_6_1/GATE.n204 VSS 0.19fF $ **FLOATING
C420 sky130_asc_pfet_01v8_lvt_6_1/GATE.n205 VSS 0.14fF $ **FLOATING
C421 porst.t7 VSS 1.97fF
C422 porst.n0 VSS 0.31fF $ **FLOATING
C423 porst.n1 VSS 0.13fF $ **FLOATING
C424 porst.t2 VSS 1.94fF
C425 porst.n2 VSS 0.53fF $ **FLOATING
C426 porst.n3 VSS 0.15fF $ **FLOATING
C427 porst.t3 VSS 1.94fF
C428 porst.n4 VSS 0.55fF $ **FLOATING
C429 porst.n5 VSS 0.15fF $ **FLOATING
C430 porst.t6 VSS 1.94fF
C431 porst.n6 VSS 0.54fF $ **FLOATING
C432 porst.n7 VSS 0.15fF $ **FLOATING
C433 porst.t1 VSS 1.94fF
C434 porst.n8 VSS 0.43fF $ **FLOATING
C435 porst.n9 VSS 0.10fF $ **FLOATING
C436 porst.n10 VSS 0.15fF $ **FLOATING
C437 porst.n11 VSS 0.10fF $ **FLOATING
C438 porst.n12 VSS 0.15fF $ **FLOATING
C439 porst.t8 VSS 1.94fF
C440 porst.n13 VSS 0.43fF $ **FLOATING
C441 porst.n14 VSS 0.10fF $ **FLOATING
C442 porst.n15 VSS 0.15fF $ **FLOATING
C443 porst.t5 VSS 1.94fF
C444 porst.n16 VSS 0.43fF $ **FLOATING
C445 porst.n17 VSS 0.10fF $ **FLOATING
C446 porst.n18 VSS 0.15fF $ **FLOATING
C447 porst.t4 VSS 1.94fF
C448 porst.n19 VSS 0.43fF $ **FLOATING
C449 porst.n20 VSS 0.10fF $ **FLOATING
C450 porst.n21 VSS 0.15fF $ **FLOATING
C451 porst.t0 VSS 1.94fF
C452 porst.n22 VSS 0.50fF $ **FLOATING
C453 porst.n23 VSS 2.36fF $ **FLOATING
C454 va.t2 VSS 1.24fF
C455 va.n0 VSS 0.34fF $ **FLOATING
C456 va.t3 VSS 1.24fF
C457 va.n1 VSS 0.35fF $ **FLOATING
C458 va.t6 VSS 1.24fF
C459 va.n2 VSS 0.34fF $ **FLOATING
C460 va.n3 VSS 0.25fF $ **FLOATING
C461 va.n4 VSS 0.56fF $ **FLOATING
C462 va.n5 VSS 0.10fF $ **FLOATING
C463 va.n6 VSS 0.10fF $ **FLOATING
C464 va.n7 VSS 0.10fF $ **FLOATING
C465 va.n8 VSS 0.52fF $ **FLOATING
C466 va.n9 VSS 0.02fF $ **FLOATING
C467 va.n10 VSS 40.66fF $ **FLOATING
C468 va.n11 VSS 13.87fF $ **FLOATING
C469 va.n12 VSS 12.41fF $ **FLOATING
C470 va.n13 VSS 13.36fF $ **FLOATING
C471 va.n14 VSS 0.13fF $ **FLOATING
C472 va.n15 VSS 0.01fF $ **FLOATING
C473 va.n16 VSS 0.00fF $ **FLOATING
C474 va.n17 VSS 0.02fF $ **FLOATING
C475 va.n18 VSS 0.00fF $ **FLOATING
C476 va.n19 VSS 0.00fF $ **FLOATING
C477 va.n20 VSS 0.00fF $ **FLOATING
C478 va.n21 VSS 0.01fF $ **FLOATING
C479 va.n22 VSS 0.00fF $ **FLOATING
C480 va.n23 VSS 0.00fF $ **FLOATING
C481 va.n24 VSS 0.01fF $ **FLOATING
C482 va.n25 VSS 0.00fF $ **FLOATING
C483 va.n26 VSS 0.01fF $ **FLOATING
C484 va.n27 VSS 0.00fF $ **FLOATING
C485 va.n28 VSS 0.01fF $ **FLOATING
C486 va.n29 VSS 0.00fF $ **FLOATING
C487 va.n30 VSS 0.00fF $ **FLOATING
C488 va.n31 VSS 0.00fF $ **FLOATING
C489 va.n32 VSS 0.01fF $ **FLOATING
C490 va.n33 VSS 0.00fF $ **FLOATING
C491 va.n34 VSS 0.00fF $ **FLOATING
C492 va.n35 VSS 0.01fF $ **FLOATING
C493 va.n36 VSS 0.00fF $ **FLOATING
C494 va.n37 VSS 0.01fF $ **FLOATING
C495 va.n38 VSS 0.00fF $ **FLOATING
C496 va.n39 VSS 0.01fF $ **FLOATING
C497 va.n40 VSS 0.00fF $ **FLOATING
C498 va.n41 VSS 0.00fF $ **FLOATING
C499 va.n42 VSS 0.00fF $ **FLOATING
C500 va.n43 VSS 0.01fF $ **FLOATING
C501 va.n44 VSS 0.00fF $ **FLOATING
C502 va.n45 VSS 0.00fF $ **FLOATING
C503 va.n46 VSS 0.01fF $ **FLOATING
C504 va.n47 VSS 0.00fF $ **FLOATING
C505 va.n48 VSS 0.01fF $ **FLOATING
C506 va.n49 VSS 0.00fF $ **FLOATING
C507 va.n50 VSS 0.01fF $ **FLOATING
C508 va.n51 VSS 0.00fF $ **FLOATING
C509 va.n52 VSS 0.00fF $ **FLOATING
C510 va.n53 VSS 0.00fF $ **FLOATING
C511 va.n54 VSS 0.01fF $ **FLOATING
C512 va.n55 VSS 0.00fF $ **FLOATING
C513 va.n56 VSS 0.00fF $ **FLOATING
C514 va.n57 VSS 0.01fF $ **FLOATING
C515 va.n58 VSS 0.00fF $ **FLOATING
C516 va.n59 VSS 0.01fF $ **FLOATING
C517 va.n60 VSS 0.00fF $ **FLOATING
C518 va.n61 VSS 0.01fF $ **FLOATING
C519 va.n62 VSS 0.00fF $ **FLOATING
C520 va.n63 VSS 0.00fF $ **FLOATING
C521 va.n64 VSS 0.00fF $ **FLOATING
C522 va.n65 VSS 0.01fF $ **FLOATING
C523 va.n66 VSS 0.00fF $ **FLOATING
C524 va.n67 VSS 0.00fF $ **FLOATING
C525 va.n68 VSS 0.01fF $ **FLOATING
C526 va.n69 VSS 0.00fF $ **FLOATING
C527 va.n70 VSS 0.01fF $ **FLOATING
C528 va.n71 VSS 0.00fF $ **FLOATING
C529 va.n72 VSS 0.01fF $ **FLOATING
C530 va.n73 VSS 0.00fF $ **FLOATING
C531 va.n74 VSS 0.00fF $ **FLOATING
C532 va.n75 VSS 0.00fF $ **FLOATING
C533 va.n76 VSS 0.01fF $ **FLOATING
C534 va.n77 VSS 0.00fF $ **FLOATING
C535 va.n78 VSS 0.00fF $ **FLOATING
C536 va.n79 VSS 0.01fF $ **FLOATING
C537 va.n80 VSS 0.00fF $ **FLOATING
C538 va.n81 VSS 0.01fF $ **FLOATING
C539 va.n82 VSS 0.00fF $ **FLOATING
C540 va.n83 VSS 0.01fF $ **FLOATING
C541 va.n84 VSS 0.00fF $ **FLOATING
C542 va.n85 VSS 0.00fF $ **FLOATING
C543 va.n86 VSS 0.00fF $ **FLOATING
C544 va.n87 VSS 0.01fF $ **FLOATING
C545 va.n88 VSS 0.00fF $ **FLOATING
C546 va.n89 VSS 0.00fF $ **FLOATING
C547 va.n90 VSS 0.01fF $ **FLOATING
C548 va.n91 VSS 0.00fF $ **FLOATING
C549 va.n92 VSS 0.01fF $ **FLOATING
C550 va.n93 VSS 0.00fF $ **FLOATING
C551 va.n94 VSS 0.01fF $ **FLOATING
C552 va.n95 VSS 0.00fF $ **FLOATING
C553 va.n96 VSS 0.00fF $ **FLOATING
C554 va.n97 VSS 0.00fF $ **FLOATING
C555 va.n98 VSS 0.01fF $ **FLOATING
C556 va.n99 VSS 0.00fF $ **FLOATING
C557 va.n100 VSS 0.00fF $ **FLOATING
C558 va.n101 VSS 0.01fF $ **FLOATING
C559 va.n102 VSS 0.00fF $ **FLOATING
C560 va.n103 VSS 0.00fF $ **FLOATING
C561 va.n104 VSS 0.00fF $ **FLOATING
C562 va.n105 VSS 0.00fF $ **FLOATING
C563 va.n106 VSS 0.01fF $ **FLOATING
C564 va.n107 VSS 0.00fF $ **FLOATING
C565 va.n108 VSS 0.01fF $ **FLOATING
C566 va.n109 VSS 0.01fF $ **FLOATING
C567 va.n110 VSS 0.00fF $ **FLOATING
C568 va.n111 VSS 0.01fF $ **FLOATING
C569 va.n112 VSS 0.00fF $ **FLOATING
C570 va.n113 VSS 0.01fF $ **FLOATING
C571 va.n114 VSS 0.00fF $ **FLOATING
C572 va.n115 VSS 0.00fF $ **FLOATING
C573 va.n116 VSS 0.00fF $ **FLOATING
C574 va.n117 VSS 0.00fF $ **FLOATING
C575 va.n118 VSS 0.01fF $ **FLOATING
C576 va.n119 VSS 0.00fF $ **FLOATING
C577 va.n120 VSS 0.01fF $ **FLOATING
C578 va.n121 VSS 0.00fF $ **FLOATING
C579 va.n122 VSS 0.01fF $ **FLOATING
C580 va.n123 VSS 0.00fF $ **FLOATING
C581 va.n124 VSS 0.01fF $ **FLOATING
C582 va.n125 VSS 0.00fF $ **FLOATING
C583 va.n126 VSS 0.00fF $ **FLOATING
C584 va.n127 VSS 0.00fF $ **FLOATING
C585 va.n128 VSS 0.00fF $ **FLOATING
C586 va.n129 VSS 0.01fF $ **FLOATING
C587 va.n130 VSS 0.00fF $ **FLOATING
C588 va.n131 VSS 0.01fF $ **FLOATING
C589 va.n132 VSS 0.00fF $ **FLOATING
C590 va.n133 VSS 0.01fF $ **FLOATING
C591 va.n134 VSS 0.00fF $ **FLOATING
C592 va.n135 VSS 0.01fF $ **FLOATING
C593 va.n136 VSS 0.00fF $ **FLOATING
C594 va.n137 VSS 0.00fF $ **FLOATING
C595 va.n138 VSS 0.00fF $ **FLOATING
C596 va.n139 VSS 0.00fF $ **FLOATING
C597 va.n140 VSS 0.01fF $ **FLOATING
C598 va.n141 VSS 0.00fF $ **FLOATING
C599 va.n142 VSS 0.01fF $ **FLOATING
C600 va.n143 VSS 0.00fF $ **FLOATING
C601 va.n144 VSS 0.01fF $ **FLOATING
C602 va.n145 VSS 0.00fF $ **FLOATING
C603 va.n146 VSS 0.01fF $ **FLOATING
C604 va.n147 VSS 0.00fF $ **FLOATING
C605 va.n148 VSS 0.00fF $ **FLOATING
C606 va.n149 VSS 0.00fF $ **FLOATING
C607 va.n150 VSS 0.00fF $ **FLOATING
C608 va.n151 VSS 0.01fF $ **FLOATING
C609 va.n152 VSS 0.00fF $ **FLOATING
C610 va.n153 VSS 0.01fF $ **FLOATING
C611 va.n154 VSS 0.00fF $ **FLOATING
C612 va.n155 VSS 0.01fF $ **FLOATING
C613 va.n156 VSS 0.00fF $ **FLOATING
C614 va.n157 VSS 0.01fF $ **FLOATING
C615 va.n158 VSS 0.00fF $ **FLOATING
C616 va.n159 VSS 0.00fF $ **FLOATING
C617 va.n160 VSS 0.00fF $ **FLOATING
C618 va.n161 VSS 0.00fF $ **FLOATING
C619 va.n162 VSS 0.01fF $ **FLOATING
C620 va.n163 VSS 0.00fF $ **FLOATING
C621 va.n164 VSS 0.01fF $ **FLOATING
C622 va.n165 VSS 0.00fF $ **FLOATING
C623 va.n166 VSS 0.01fF $ **FLOATING
C624 va.n167 VSS 0.00fF $ **FLOATING
C625 va.n168 VSS 0.01fF $ **FLOATING
C626 va.n169 VSS 0.00fF $ **FLOATING
C627 va.n170 VSS 0.00fF $ **FLOATING
C628 va.n171 VSS 0.00fF $ **FLOATING
C629 va.n172 VSS 0.00fF $ **FLOATING
C630 va.n173 VSS 0.01fF $ **FLOATING
C631 va.n174 VSS 0.00fF $ **FLOATING
C632 va.n175 VSS 0.01fF $ **FLOATING
C633 va.n176 VSS 0.00fF $ **FLOATING
C634 va.n177 VSS 0.01fF $ **FLOATING
C635 va.n178 VSS 0.00fF $ **FLOATING
C636 va.n179 VSS 0.01fF $ **FLOATING
C637 va.n180 VSS 0.00fF $ **FLOATING
C638 va.n181 VSS 0.00fF $ **FLOATING
C639 va.n182 VSS 0.00fF $ **FLOATING
C640 va.n183 VSS 0.00fF $ **FLOATING
C641 va.n184 VSS 0.01fF $ **FLOATING
C642 va.n185 VSS 0.00fF $ **FLOATING
C643 va.n186 VSS 0.01fF $ **FLOATING
C644 va.n187 VSS 0.00fF $ **FLOATING
C645 va.n188 VSS 0.01fF $ **FLOATING
C646 va.n189 VSS 0.01fF $ **FLOATING
C647 va.n190 VSS 0.00fF $ **FLOATING
C648 va.n191 VSS 0.02fF $ **FLOATING
C649 va.n192 VSS 0.10fF $ **FLOATING
C650 va.n193 VSS 27.18fF $ **FLOATING
C651 va.n194 VSS 26.34fF $ **FLOATING
C652 va.n195 VSS 2.99fF $ **FLOATING
C653 va.n196 VSS 29.80fF $ **FLOATING
C654 va.n197 VSS 0.58fF $ **FLOATING
C655 va.n198 VSS 0.02fF $ **FLOATING
C656 va.n199 VSS 0.11fF $ **FLOATING
C657 va.n200 VSS 0.11fF $ **FLOATING
C658 va.n201 VSS 0.22fF $ **FLOATING
C659 va.n202 VSS 0.11fF $ **FLOATING
C660 va.n203 VSS 0.02fF $ **FLOATING
C661 va.n204 VSS 0.12fF $ **FLOATING
C662 va.n205 VSS 0.04fF $ **FLOATING
C663 va.n206 VSS 0.02fF $ **FLOATING
C664 va.n207 VSS 0.03fF $ **FLOATING
C665 va.n208 VSS 0.06fF $ **FLOATING
C666 va.n209 VSS 0.09fF $ **FLOATING
C667 va.n210 VSS 0.02fF $ **FLOATING
C668 va.n211 VSS 0.14fF $ **FLOATING
C669 va.n212 VSS 0.02fF $ **FLOATING
C670 va.n213 VSS 0.12fF $ **FLOATING
C671 va.n214 VSS 0.03fF $ **FLOATING
C672 va.n215 VSS 0.02fF $ **FLOATING
C673 va.n216 VSS 0.02fF $ **FLOATING
C674 va.n217 VSS 0.10fF $ **FLOATING
C675 va.n218 VSS 0.11fF $ **FLOATING
C676 va.n219 VSS 0.14fF $ **FLOATING
C677 va.n220 VSS 0.24fF $ **FLOATING
C678 va.n221 VSS 0.14fF $ **FLOATING
C679 va.n222 VSS 0.14fF $ **FLOATING
C680 va.n223 VSS 0.12fF $ **FLOATING
C681 va.n224 VSS 0.24fF $ **FLOATING
C682 va.n225 VSS 0.14fF $ **FLOATING
C683 va.n226 VSS 0.12fF $ **FLOATING
C684 va.n227 VSS 0.23fF $ **FLOATING
C685 va.n228 VSS 0.14fF $ **FLOATING
C686 va.n229 VSS 0.27fF $ **FLOATING
C687 va.t0 VSS 1.24fF
C688 va.n230 VSS 0.30fF $ **FLOATING
C689 va.n231 VSS 0.15fF $ **FLOATING
C690 va.n232 VSS 0.07fF $ **FLOATING
C691 va.n233 VSS 0.10fF $ **FLOATING
C692 va.t4 VSS 1.24fF
C693 va.n234 VSS 0.28fF $ **FLOATING
C694 va.n235 VSS 0.07fF $ **FLOATING
C695 va.n236 VSS 0.09fF $ **FLOATING
C696 va.t5 VSS 1.24fF
C697 va.n237 VSS 0.28fF $ **FLOATING
C698 va.n238 VSS 0.07fF $ **FLOATING
C699 va.n239 VSS 0.09fF $ **FLOATING
C700 va.t8 VSS 1.24fF
C701 va.n240 VSS 0.28fF $ **FLOATING
C702 va.n241 VSS 0.07fF $ **FLOATING
C703 va.n242 VSS 0.09fF $ **FLOATING
C704 va.t1 VSS 1.24fF
C705 va.n243 VSS 0.28fF $ **FLOATING
C706 va.n244 VSS 0.07fF $ **FLOATING
C707 va.n245 VSS 0.09fF $ **FLOATING
C708 va.n246 VSS 0.09fF $ **FLOATING
C709 va.n247 VSS 0.09fF $ **FLOATING
C710 va.n248 VSS 0.09fF $ **FLOATING
C711 va.t7 VSS 1.26fF
C712 va.n249 VSS 0.20fF $ **FLOATING
C713 va.n250 VSS 0.08fF $ **FLOATING
C714 vb.t7 VSS 1.78fF
C715 vb.n0 VSS 0.28fF $ **FLOATING
C716 vb.t2 VSS 1.75fF
C717 vb.n1 VSS 0.48fF $ **FLOATING
C718 vb.t3 VSS 1.75fF
C719 vb.n2 VSS 0.50fF $ **FLOATING
C720 vb.t6 VSS 1.75fF
C721 vb.n3 VSS 0.48fF $ **FLOATING
C722 vb.n4 VSS 2.12fF $ **FLOATING
C723 vb.n5 VSS 1.12fF $ **FLOATING
C724 vb.n6 VSS 0.03fF $ **FLOATING
C725 vb.n7 VSS 0.01fF $ **FLOATING
C726 vb.n8 VSS 0.01fF $ **FLOATING
C727 vb.n9 VSS 0.00fF $ **FLOATING
C728 vb.n10 VSS 0.00fF $ **FLOATING
C729 vb.n11 VSS 0.00fF $ **FLOATING
C730 vb.n12 VSS 0.01fF $ **FLOATING
C731 vb.n13 VSS 0.00fF $ **FLOATING
C732 vb.n14 VSS 0.00fF $ **FLOATING
C733 vb.n15 VSS 0.01fF $ **FLOATING
C734 vb.n16 VSS 0.00fF $ **FLOATING
C735 vb.n17 VSS 0.01fF $ **FLOATING
C736 vb.n18 VSS 0.00fF $ **FLOATING
C737 vb.n19 VSS 0.01fF $ **FLOATING
C738 vb.n20 VSS 0.00fF $ **FLOATING
C739 vb.n21 VSS 0.00fF $ **FLOATING
C740 vb.n22 VSS 0.00fF $ **FLOATING
C741 vb.n23 VSS 0.01fF $ **FLOATING
C742 vb.n24 VSS 0.00fF $ **FLOATING
C743 vb.n25 VSS 0.00fF $ **FLOATING
C744 vb.n26 VSS 0.01fF $ **FLOATING
C745 vb.n27 VSS 0.00fF $ **FLOATING
C746 vb.n28 VSS 0.01fF $ **FLOATING
C747 vb.n29 VSS 0.00fF $ **FLOATING
C748 vb.n30 VSS 0.01fF $ **FLOATING
C749 vb.n31 VSS 0.00fF $ **FLOATING
C750 vb.n32 VSS 0.00fF $ **FLOATING
C751 vb.n33 VSS 0.00fF $ **FLOATING
C752 vb.n34 VSS 0.01fF $ **FLOATING
C753 vb.n35 VSS 0.00fF $ **FLOATING
C754 vb.n36 VSS 0.00fF $ **FLOATING
C755 vb.n37 VSS 0.01fF $ **FLOATING
C756 vb.n38 VSS 0.00fF $ **FLOATING
C757 vb.n39 VSS 0.01fF $ **FLOATING
C758 vb.n40 VSS 0.00fF $ **FLOATING
C759 vb.n41 VSS 0.01fF $ **FLOATING
C760 vb.n42 VSS 0.00fF $ **FLOATING
C761 vb.n43 VSS 0.00fF $ **FLOATING
C762 vb.n44 VSS 0.00fF $ **FLOATING
C763 vb.n45 VSS 0.01fF $ **FLOATING
C764 vb.n46 VSS 0.00fF $ **FLOATING
C765 vb.n47 VSS 0.00fF $ **FLOATING
C766 vb.n48 VSS 0.01fF $ **FLOATING
C767 vb.n49 VSS 0.00fF $ **FLOATING
C768 vb.n50 VSS 0.01fF $ **FLOATING
C769 vb.n51 VSS 0.00fF $ **FLOATING
C770 vb.n52 VSS 0.01fF $ **FLOATING
C771 vb.n53 VSS 0.00fF $ **FLOATING
C772 vb.n54 VSS 0.00fF $ **FLOATING
C773 vb.n55 VSS 0.00fF $ **FLOATING
C774 vb.n56 VSS 0.01fF $ **FLOATING
C775 vb.n57 VSS 0.00fF $ **FLOATING
C776 vb.n58 VSS 0.00fF $ **FLOATING
C777 vb.n59 VSS 0.01fF $ **FLOATING
C778 vb.n60 VSS 0.00fF $ **FLOATING
C779 vb.n61 VSS 0.01fF $ **FLOATING
C780 vb.n62 VSS 0.00fF $ **FLOATING
C781 vb.n63 VSS 0.01fF $ **FLOATING
C782 vb.n64 VSS 0.00fF $ **FLOATING
C783 vb.n65 VSS 0.00fF $ **FLOATING
C784 vb.n66 VSS 0.00fF $ **FLOATING
C785 vb.n67 VSS 0.01fF $ **FLOATING
C786 vb.n68 VSS 0.00fF $ **FLOATING
C787 vb.n69 VSS 0.00fF $ **FLOATING
C788 vb.n70 VSS 0.01fF $ **FLOATING
C789 vb.n71 VSS 0.00fF $ **FLOATING
C790 vb.n72 VSS 0.01fF $ **FLOATING
C791 vb.n73 VSS 0.00fF $ **FLOATING
C792 vb.n74 VSS 0.01fF $ **FLOATING
C793 vb.n75 VSS 0.00fF $ **FLOATING
C794 vb.n76 VSS 0.00fF $ **FLOATING
C795 vb.n77 VSS 0.00fF $ **FLOATING
C796 vb.n78 VSS 0.01fF $ **FLOATING
C797 vb.n79 VSS 0.00fF $ **FLOATING
C798 vb.n80 VSS 0.00fF $ **FLOATING
C799 vb.n81 VSS 0.01fF $ **FLOATING
C800 vb.n82 VSS 0.00fF $ **FLOATING
C801 vb.n83 VSS 0.01fF $ **FLOATING
C802 vb.n84 VSS 0.00fF $ **FLOATING
C803 vb.n85 VSS 0.01fF $ **FLOATING
C804 vb.n86 VSS 0.00fF $ **FLOATING
C805 vb.n87 VSS 0.00fF $ **FLOATING
C806 vb.n88 VSS 0.00fF $ **FLOATING
C807 vb.n89 VSS 0.01fF $ **FLOATING
C808 vb.n90 VSS 0.01fF $ **FLOATING
C809 vb.n91 VSS 0.00fF $ **FLOATING
C810 vb.n92 VSS 0.01fF $ **FLOATING
C811 vb.n93 VSS 0.00fF $ **FLOATING
C812 vb.n94 VSS 0.00fF $ **FLOATING
C813 vb.n95 VSS 0.00fF $ **FLOATING
C814 vb.n96 VSS 0.00fF $ **FLOATING
C815 vb.n97 VSS 0.02fF $ **FLOATING
C816 vb.n98 VSS 0.01fF $ **FLOATING
C817 vb.n99 VSS 0.00fF $ **FLOATING
C818 vb.n100 VSS 0.01fF $ **FLOATING
C819 vb.n101 VSS 0.00fF $ **FLOATING
C820 vb.n102 VSS 0.01fF $ **FLOATING
C821 vb.n103 VSS 0.00fF $ **FLOATING
C822 vb.n104 VSS 0.01fF $ **FLOATING
C823 vb.n105 VSS 0.00fF $ **FLOATING
C824 vb.n106 VSS 0.00fF $ **FLOATING
C825 vb.n107 VSS 0.00fF $ **FLOATING
C826 vb.n108 VSS 0.00fF $ **FLOATING
C827 vb.n109 VSS 0.01fF $ **FLOATING
C828 vb.n110 VSS 0.00fF $ **FLOATING
C829 vb.n111 VSS 0.01fF $ **FLOATING
C830 vb.n112 VSS 0.00fF $ **FLOATING
C831 vb.n113 VSS 0.01fF $ **FLOATING
C832 vb.n114 VSS 0.00fF $ **FLOATING
C833 vb.n115 VSS 0.01fF $ **FLOATING
C834 vb.n116 VSS 0.00fF $ **FLOATING
C835 vb.n117 VSS 0.00fF $ **FLOATING
C836 vb.n118 VSS 0.00fF $ **FLOATING
C837 vb.n119 VSS 0.00fF $ **FLOATING
C838 vb.n120 VSS 0.01fF $ **FLOATING
C839 vb.n121 VSS 0.00fF $ **FLOATING
C840 vb.n122 VSS 0.01fF $ **FLOATING
C841 vb.n123 VSS 0.00fF $ **FLOATING
C842 vb.n124 VSS 0.01fF $ **FLOATING
C843 vb.n125 VSS 0.00fF $ **FLOATING
C844 vb.n126 VSS 0.01fF $ **FLOATING
C845 vb.n127 VSS 0.00fF $ **FLOATING
C846 vb.n128 VSS 0.00fF $ **FLOATING
C847 vb.n129 VSS 0.00fF $ **FLOATING
C848 vb.n130 VSS 0.00fF $ **FLOATING
C849 vb.n131 VSS 0.01fF $ **FLOATING
C850 vb.n132 VSS 0.00fF $ **FLOATING
C851 vb.n133 VSS 0.01fF $ **FLOATING
C852 vb.n134 VSS 0.00fF $ **FLOATING
C853 vb.n135 VSS 0.01fF $ **FLOATING
C854 vb.n136 VSS 0.00fF $ **FLOATING
C855 vb.n137 VSS 0.01fF $ **FLOATING
C856 vb.n138 VSS 0.00fF $ **FLOATING
C857 vb.n139 VSS 0.00fF $ **FLOATING
C858 vb.n140 VSS 0.00fF $ **FLOATING
C859 vb.n141 VSS 0.00fF $ **FLOATING
C860 vb.n142 VSS 0.01fF $ **FLOATING
C861 vb.n143 VSS 0.00fF $ **FLOATING
C862 vb.n144 VSS 0.01fF $ **FLOATING
C863 vb.n145 VSS 0.00fF $ **FLOATING
C864 vb.n146 VSS 0.01fF $ **FLOATING
C865 vb.n147 VSS 0.00fF $ **FLOATING
C866 vb.n148 VSS 0.01fF $ **FLOATING
C867 vb.n149 VSS 0.00fF $ **FLOATING
C868 vb.n150 VSS 0.00fF $ **FLOATING
C869 vb.n151 VSS 0.00fF $ **FLOATING
C870 vb.n152 VSS 0.00fF $ **FLOATING
C871 vb.n153 VSS 0.01fF $ **FLOATING
C872 vb.n154 VSS 0.00fF $ **FLOATING
C873 vb.n155 VSS 0.01fF $ **FLOATING
C874 vb.n156 VSS 0.00fF $ **FLOATING
C875 vb.n157 VSS 0.01fF $ **FLOATING
C876 vb.n158 VSS 0.00fF $ **FLOATING
C877 vb.n159 VSS 0.01fF $ **FLOATING
C878 vb.n160 VSS 0.00fF $ **FLOATING
C879 vb.n161 VSS 0.00fF $ **FLOATING
C880 vb.n162 VSS 0.00fF $ **FLOATING
C881 vb.n163 VSS 0.00fF $ **FLOATING
C882 vb.n164 VSS 0.01fF $ **FLOATING
C883 vb.n165 VSS 0.00fF $ **FLOATING
C884 vb.n166 VSS 0.01fF $ **FLOATING
C885 vb.n167 VSS 0.00fF $ **FLOATING
C886 vb.n168 VSS 0.01fF $ **FLOATING
C887 vb.n169 VSS 0.00fF $ **FLOATING
C888 vb.n170 VSS 0.01fF $ **FLOATING
C889 vb.n171 VSS 0.00fF $ **FLOATING
C890 vb.n172 VSS 0.00fF $ **FLOATING
C891 vb.n173 VSS 0.02fF $ **FLOATING
C892 vb.n174 VSS 0.01fF $ **FLOATING
C893 vb.n175 VSS 0.03fF $ **FLOATING
C894 vb.n176 VSS 0.04fF $ **FLOATING
C895 vb.n177 VSS 10.08fF $ **FLOATING
C896 vb.n178 VSS 30.50fF $ **FLOATING
C897 vb.t0 VSS 1.75fF
C898 vb.n179 VSS 0.45fF $ **FLOATING
C899 vb.n180 VSS 0.30fF $ **FLOATING
C900 vb.n181 VSS 0.09fF $ **FLOATING
C901 vb.n182 VSS 0.13fF $ **FLOATING
C902 vb.t4 VSS 1.75fF
C903 vb.n183 VSS 0.39fF $ **FLOATING
C904 vb.n184 VSS 0.09fF $ **FLOATING
C905 vb.n185 VSS 0.13fF $ **FLOATING
C906 vb.t5 VSS 1.75fF
C907 vb.n186 VSS 0.39fF $ **FLOATING
C908 vb.n187 VSS 0.09fF $ **FLOATING
C909 vb.n188 VSS 0.13fF $ **FLOATING
C910 vb.t8 VSS 1.75fF
C911 vb.n189 VSS 0.39fF $ **FLOATING
C912 vb.n190 VSS 0.09fF $ **FLOATING
C913 vb.n191 VSS 0.13fF $ **FLOATING
C914 vb.t1 VSS 1.75fF
C915 vb.n192 VSS 0.39fF $ **FLOATING
C916 vb.n193 VSS 0.09fF $ **FLOATING
C917 vb.n194 VSS 0.13fF $ **FLOATING
C918 vb.n195 VSS 0.13fF $ **FLOATING
C919 vb.n196 VSS 0.13fF $ **FLOATING
C920 vb.n197 VSS 0.13fF $ **FLOATING
C921 vb.n198 VSS 0.12fF $ **FLOATING
C922  VSS 31.69fF $ **FLOATING
C923 VDD.n0 VSS 61.55fF $ **FLOATING
C924 VDD.n3 VSS 0.01fF $ **FLOATING
C925 VDD.n4 VSS 0.07fF $ **FLOATING
C926 VDD.n6 VSS 0.01fF $ **FLOATING
C927 VDD.n7 VSS 0.00fF $ **FLOATING
C928 VDD.n8 VSS 0.01fF $ **FLOATING
C929 VDD.n9 VSS 0.01fF $ **FLOATING
C930 VDD.n10 VSS 0.03fF $ **FLOATING
C931 VDD.n11 VSS 0.09fF $ **FLOATING
C932 VDD.n12 VSS 0.01fF $ **FLOATING
C933 VDD.n13 VSS 0.07fF $ **FLOATING
C934 VDD.n14 VSS 0.00fF $ **FLOATING
C935 VDD.n15 VSS 0.01fF $ **FLOATING
C936 VDD.n16 VSS 0.03fF $ **FLOATING
C937 VDD.n17 VSS 0.04fF $ **FLOATING
C938 VDD.n18 VSS 0.03fF $ **FLOATING
C939 VDD.n19 VSS 0.04fF $ **FLOATING
C940 VDD.n20 VSS 0.00fF $ **FLOATING
C941 VDD.n21 VSS 0.07fF $ **FLOATING
C942 VDD.n22 VSS 0.00fF $ **FLOATING
C943 VDD.n24 VSS 0.01fF $ **FLOATING
C944 VDD.n25 VSS 0.07fF $ **FLOATING
C945 VDD.n27 VSS 0.01fF $ **FLOATING
C946 VDD.n28 VSS 0.00fF $ **FLOATING
C947 VDD.n29 VSS 0.01fF $ **FLOATING
C948 VDD.n30 VSS 0.01fF $ **FLOATING
C949 VDD.n31 VSS 0.03fF $ **FLOATING
C950 VDD.n32 VSS 0.09fF $ **FLOATING
C951 VDD.n33 VSS 0.01fF $ **FLOATING
C952 VDD.n34 VSS 0.07fF $ **FLOATING
C953 VDD.n35 VSS 0.00fF $ **FLOATING
C954 VDD.n36 VSS 0.01fF $ **FLOATING
C955 VDD.n37 VSS 0.03fF $ **FLOATING
C956 VDD.n38 VSS 0.04fF $ **FLOATING
C957 VDD.n39 VSS 0.03fF $ **FLOATING
C958 VDD.n40 VSS 0.04fF $ **FLOATING
C959 VDD.n41 VSS 0.00fF $ **FLOATING
C960 VDD.n42 VSS 0.07fF $ **FLOATING
C961 VDD.n43 VSS 0.00fF $ **FLOATING
C962 VDD.n45 VSS 0.01fF $ **FLOATING
C963 VDD.n46 VSS 0.07fF $ **FLOATING
C964 VDD.n48 VSS 0.01fF $ **FLOATING
C965 VDD.n49 VSS 0.00fF $ **FLOATING
C966 VDD.n50 VSS 0.01fF $ **FLOATING
C967 VDD.n51 VSS 0.01fF $ **FLOATING
C968 VDD.n52 VSS 0.03fF $ **FLOATING
C969 VDD.n53 VSS 0.09fF $ **FLOATING
C970 VDD.n54 VSS 0.01fF $ **FLOATING
C971 VDD.n55 VSS 0.07fF $ **FLOATING
C972 VDD.n56 VSS 0.00fF $ **FLOATING
C973 VDD.n57 VSS 0.01fF $ **FLOATING
C974 VDD.n58 VSS 0.03fF $ **FLOATING
C975 VDD.n59 VSS 0.04fF $ **FLOATING
C976 VDD.n60 VSS 0.03fF $ **FLOATING
C977 VDD.n61 VSS 0.04fF $ **FLOATING
C978 VDD.n62 VSS 0.00fF $ **FLOATING
C979 VDD.n63 VSS 0.07fF $ **FLOATING
C980 VDD.n64 VSS 0.00fF $ **FLOATING
C981 VDD.n66 VSS 0.01fF $ **FLOATING
C982 VDD.n67 VSS 0.07fF $ **FLOATING
C983 VDD.n69 VSS 0.01fF $ **FLOATING
C984 VDD.n70 VSS 0.00fF $ **FLOATING
C985 VDD.n71 VSS 0.01fF $ **FLOATING
C986 VDD.n72 VSS 0.01fF $ **FLOATING
C987 VDD.n73 VSS 0.03fF $ **FLOATING
C988 VDD.n74 VSS 0.09fF $ **FLOATING
C989 VDD.n75 VSS 0.01fF $ **FLOATING
C990 VDD.n76 VSS 0.07fF $ **FLOATING
C991 VDD.n77 VSS 0.00fF $ **FLOATING
C992 VDD.n78 VSS 0.01fF $ **FLOATING
C993 VDD.n79 VSS 0.03fF $ **FLOATING
C994 VDD.n80 VSS 0.04fF $ **FLOATING
C995 VDD.n81 VSS 0.03fF $ **FLOATING
C996 VDD.n82 VSS 0.04fF $ **FLOATING
C997 VDD.n83 VSS 0.00fF $ **FLOATING
C998 VDD.n84 VSS 0.07fF $ **FLOATING
C999 VDD.n85 VSS 0.00fF $ **FLOATING
C1000 VDD.n87 VSS 0.01fF $ **FLOATING
C1001 VDD.n88 VSS 0.07fF $ **FLOATING
C1002 VDD.n90 VSS 0.01fF $ **FLOATING
C1003 VDD.n91 VSS 0.00fF $ **FLOATING
C1004 VDD.n92 VSS 0.01fF $ **FLOATING
C1005 VDD.n93 VSS 0.01fF $ **FLOATING
C1006 VDD.n94 VSS 0.03fF $ **FLOATING
C1007 VDD.n95 VSS 0.09fF $ **FLOATING
C1008 VDD.n96 VSS 0.01fF $ **FLOATING
C1009 VDD.n97 VSS 0.07fF $ **FLOATING
C1010 VDD.n98 VSS 0.00fF $ **FLOATING
C1011 VDD.n99 VSS 0.01fF $ **FLOATING
C1012 VDD.n100 VSS 0.03fF $ **FLOATING
C1013 VDD.n101 VSS 0.04fF $ **FLOATING
C1014 VDD.n102 VSS 0.03fF $ **FLOATING
C1015 VDD.n103 VSS 0.04fF $ **FLOATING
C1016 VDD.n104 VSS 0.00fF $ **FLOATING
C1017 VDD.n105 VSS 0.07fF $ **FLOATING
C1018 VDD.n106 VSS 0.00fF $ **FLOATING
C1019 VDD.n108 VSS 0.01fF $ **FLOATING
C1020 VDD.n109 VSS 0.07fF $ **FLOATING
C1021 VDD.n111 VSS 0.01fF $ **FLOATING
C1022 VDD.n112 VSS 0.00fF $ **FLOATING
C1023 VDD.n113 VSS 0.01fF $ **FLOATING
C1024 VDD.n114 VSS 0.01fF $ **FLOATING
C1025 VDD.n115 VSS 0.03fF $ **FLOATING
C1026 VDD.n116 VSS 0.09fF $ **FLOATING
C1027 VDD.n117 VSS 0.01fF $ **FLOATING
C1028 VDD.n118 VSS 0.07fF $ **FLOATING
C1029 VDD.n119 VSS 0.00fF $ **FLOATING
C1030 VDD.n120 VSS 0.01fF $ **FLOATING
C1031 VDD.n121 VSS 0.03fF $ **FLOATING
C1032 VDD.n122 VSS 0.04fF $ **FLOATING
C1033 VDD.n123 VSS 0.03fF $ **FLOATING
C1034 VDD.n124 VSS 0.04fF $ **FLOATING
C1035 VDD.n125 VSS 0.00fF $ **FLOATING
C1036 VDD.n126 VSS 0.07fF $ **FLOATING
C1037 VDD.n127 VSS 0.00fF $ **FLOATING
C1038 VDD.n129 VSS 0.01fF $ **FLOATING
C1039 VDD.n130 VSS 0.07fF $ **FLOATING
C1040 VDD.n132 VSS 0.01fF $ **FLOATING
C1041 VDD.n133 VSS 0.00fF $ **FLOATING
C1042 VDD.n134 VSS 0.01fF $ **FLOATING
C1043 VDD.n135 VSS 0.01fF $ **FLOATING
C1044 VDD.n136 VSS 0.03fF $ **FLOATING
C1045 VDD.n137 VSS 0.09fF $ **FLOATING
C1046 VDD.n138 VSS 0.01fF $ **FLOATING
C1047 VDD.n139 VSS 0.07fF $ **FLOATING
C1048 VDD.n140 VSS 0.00fF $ **FLOATING
C1049 VDD.n141 VSS 0.01fF $ **FLOATING
C1050 VDD.n142 VSS 0.03fF $ **FLOATING
C1051 VDD.n143 VSS 0.04fF $ **FLOATING
C1052 VDD.n144 VSS 0.03fF $ **FLOATING
C1053 VDD.n145 VSS 0.04fF $ **FLOATING
C1054 VDD.n146 VSS 0.00fF $ **FLOATING
C1055 VDD.n147 VSS 0.07fF $ **FLOATING
C1056 VDD.n148 VSS 0.00fF $ **FLOATING
C1057 VDD.n150 VSS 0.01fF $ **FLOATING
C1058 VDD.n151 VSS 0.07fF $ **FLOATING
C1059 VDD.n153 VSS 0.01fF $ **FLOATING
C1060 VDD.n154 VSS 0.00fF $ **FLOATING
C1061 VDD.n155 VSS 0.01fF $ **FLOATING
C1062 VDD.n156 VSS 0.01fF $ **FLOATING
C1063 VDD.n157 VSS 0.03fF $ **FLOATING
C1064 VDD.n158 VSS 0.09fF $ **FLOATING
C1065 VDD.n159 VSS 0.01fF $ **FLOATING
C1066 VDD.n160 VSS 0.07fF $ **FLOATING
C1067 VDD.n161 VSS 0.00fF $ **FLOATING
C1068 VDD.n162 VSS 0.01fF $ **FLOATING
C1069 VDD.n163 VSS 0.03fF $ **FLOATING
C1070 VDD.n164 VSS 0.04fF $ **FLOATING
C1071 VDD.n165 VSS 0.03fF $ **FLOATING
C1072 VDD.n166 VSS 0.04fF $ **FLOATING
C1073 VDD.n167 VSS 0.00fF $ **FLOATING
C1074 VDD.n168 VSS 0.07fF $ **FLOATING
C1075 VDD.n169 VSS 0.00fF $ **FLOATING
C1076 VDD.n170 VSS 4.15fF $ **FLOATING
C1077 VDD.n172 VSS 0.03fF $ **FLOATING
C1078 VDD.n173 VSS 0.01fF $ **FLOATING
C1079 VDD.n174 VSS 0.00fF $ **FLOATING
C1080 VDD.n175 VSS 0.01fF $ **FLOATING
C1081 VDD.n176 VSS 0.01fF $ **FLOATING
C1082 VDD.n177 VSS 0.09fF $ **FLOATING
C1083 VDD.n178 VSS 0.01fF $ **FLOATING
C1084 VDD.n179 VSS 0.07fF $ **FLOATING
C1085 VDD.n180 VSS 0.01fF $ **FLOATING
C1086 VDD.n181 VSS 0.07fF $ **FLOATING
C1087 VDD.n182 VSS 0.03fF $ **FLOATING
C1088 VDD.n183 VSS 0.03fF $ **FLOATING
C1089 VDD.n184 VSS 0.03fF $ **FLOATING
C1090 VDD.n185 VSS 0.06fF $ **FLOATING
C1091 VDD.n186 VSS 0.13fF $ **FLOATING
C1092 VDD.n187 VSS 12.46fF $ **FLOATING
C1093 VDD.n188 VSS 0.70fF $ **FLOATING
C1094 VDD.n189 VSS 12.46fF $ **FLOATING
C1095 VDD.n190 VSS 0.13fF $ **FLOATING
C1096 VDD.n191 VSS 0.70fF $ **FLOATING
C1097 VDD.n192 VSS 0.07fF $ **FLOATING
C1098 VDD.n193 VSS 60.75fF $ **FLOATING
C1099 VDD.n194 VSS 61.56fF $ **FLOATING
C1100 VDD.n195 VSS 4.15fF $ **FLOATING
C1101 VDD.n197 VSS 0.03fF $ **FLOATING
C1102 VDD.n198 VSS 0.01fF $ **FLOATING
C1103 VDD.n199 VSS 0.00fF $ **FLOATING
C1104 VDD.n200 VSS 0.01fF $ **FLOATING
C1105 VDD.n201 VSS 0.01fF $ **FLOATING
C1106 VDD.n202 VSS 0.09fF $ **FLOATING
C1107 VDD.n203 VSS 0.01fF $ **FLOATING
C1108 VDD.n204 VSS 0.07fF $ **FLOATING
C1109 VDD.n205 VSS 0.01fF $ **FLOATING
C1110 VDD.n206 VSS 0.07fF $ **FLOATING
C1111 VDD.n207 VSS 0.01fF $ **FLOATING
C1112 VDD.n208 VSS 0.03fF $ **FLOATING
C1113 VDD.n209 VSS 0.01fF $ **FLOATING
C1114 VDD.n210 VSS 0.00fF $ **FLOATING
C1115 VDD.n211 VSS 0.01fF $ **FLOATING
C1116 VDD.n212 VSS 0.01fF $ **FLOATING
C1117 VDD.n213 VSS 0.09fF $ **FLOATING
C1118 VDD.n214 VSS 0.01fF $ **FLOATING
C1119 VDD.n215 VSS 0.07fF $ **FLOATING
C1120 VDD.n216 VSS 0.01fF $ **FLOATING
C1121 VDD.n217 VSS 0.07fF $ **FLOATING
C1122 VDD.n218 VSS 0.01fF $ **FLOATING
C1123 VDD.n219 VSS 0.07fF $ **FLOATING
C1124 VDD.n220 VSS 0.03fF $ **FLOATING
C1125 VDD.t14 VSS 0.05fF
C1126 VDD.t35 VSS 0.05fF
C1127 VDD.n221 VSS 0.37fF $ **FLOATING
C1128 VDD.t2 VSS 0.05fF
C1129 VDD.t17 VSS 0.05fF
C1130 VDD.n222 VSS 0.37fF $ **FLOATING
C1131 VDD.t11 VSS 0.05fF
C1132 VDD.t5 VSS 0.05fF
C1133 VDD.n223 VSS 0.37fF $ **FLOATING
C1134 VDD.t29 VSS 0.05fF
C1135 VDD.t23 VSS 0.05fF
C1136 VDD.n224 VSS 0.37fF $ **FLOATING
C1137 VDD.t20 VSS 0.05fF
C1138 VDD.t8 VSS 0.05fF
C1139 VDD.n225 VSS 0.37fF $ **FLOATING
C1140 VDD.t32 VSS 0.05fF
C1141 VDD.t26 VSS 0.05fF
C1142 VDD.n226 VSS 0.37fF $ **FLOATING
C1143 VDD.n227 VSS 0.08fF $ **FLOATING
C1144 VDD.n228 VSS 0.11fF $ **FLOATING
C1145 VDD.n229 VSS 0.11fF $ **FLOATING
C1146 VDD.n230 VSS 0.11fF $ **FLOATING
C1147 VDD.n231 VSS 0.11fF $ **FLOATING
C1148 VDD.n232 VSS 0.08fF $ **FLOATING
C1149 VDD.n233 VSS 0.13fF $ **FLOATING
C1150 VDD.n234 VSS 0.06fF $ **FLOATING
C1151 VDD.t16 VSS 1.34fF
C1152 VDD.n235 VSS 0.06fF $ **FLOATING
C1153 VDD.n236 VSS 0.13fF $ **FLOATING
C1154 VDD.n237 VSS 0.05fF $ **FLOATING
C1155 VDD.t31 VSS 2.30fF
C1156 VDD.t25 VSS 2.02fF
C1157 VDD.t19 VSS 2.02fF
C1158 VDD.t7 VSS 1.66fF
C1159 VDD.n238 VSS 0.06fF $ **FLOATING
C1160 VDD.t30 VSS 1.22fF
C1161 VDD.t18 VSS 1.22fF
C1162 VDD.n239 VSS 0.28fF $ **FLOATING
C1163 VDD.n240 VSS 0.06fF $ **FLOATING
C1164 VDD.t21 VSS 1.22fF
C1165 VDD.n241 VSS 0.32fF $ **FLOATING
C1166 VDD.t9 VSS 1.22fF
C1167 VDD.n242 VSS 0.33fF $ **FLOATING
C1168 VDD.n243 VSS 0.06fF $ **FLOATING
C1169 VDD.t15 VSS 1.22fF
C1170 VDD.n244 VSS 0.28fF $ **FLOATING
C1171 VDD.t33 VSS 1.31fF
C1172 VDD.n245 VSS 0.37fF $ **FLOATING
C1173 VDD.t12 VSS 1.22fF
C1174 VDD.n246 VSS 0.29fF $ **FLOATING
C1175 VDD.n247 VSS 0.04fF $ **FLOATING
C1176 VDD.n248 VSS 0.10fF $ **FLOATING
C1177 VDD.n249 VSS 0.06fF $ **FLOATING
C1178 VDD.n250 VSS 0.04fF $ **FLOATING
C1179 VDD.t0 VSS 1.22fF
C1180 VDD.n251 VSS 0.28fF $ **FLOATING
C1181 VDD.n252 VSS 0.04fF $ **FLOATING
C1182 VDD.t3 VSS 1.22fF
C1183 VDD.n253 VSS 0.28fF $ **FLOATING
C1184 VDD.n254 VSS 0.04fF $ **FLOATING
C1185 VDD.n255 VSS 0.06fF $ **FLOATING
C1186 VDD.n256 VSS 0.06fF $ **FLOATING
C1187 VDD.n257 VSS 0.06fF $ **FLOATING
C1188 VDD.n258 VSS 0.06fF $ **FLOATING
C1189 VDD.n259 VSS 0.04fF $ **FLOATING
C1190 VDD.t27 VSS 1.22fF
C1191 VDD.n260 VSS 0.28fF $ **FLOATING
C1192 VDD.n261 VSS 0.04fF $ **FLOATING
C1193 VDD.t6 VSS 1.22fF
C1194 VDD.n262 VSS 0.28fF $ **FLOATING
C1195 VDD.n263 VSS 0.04fF $ **FLOATING
C1196 VDD.n264 VSS 0.06fF $ **FLOATING
C1197 VDD.n265 VSS 0.06fF $ **FLOATING
C1198 VDD.n266 VSS 0.04fF $ **FLOATING
C1199 VDD.t24 VSS 1.22fF
C1200 VDD.n267 VSS 0.28fF $ **FLOATING
C1201 VDD.n268 VSS 0.04fF $ **FLOATING
C1202 VDD.n269 VSS 0.33fF $ **FLOATING
C1203 VDD.n270 VSS 0.05fF $ **FLOATING
C1204 VDD.n271 VSS 0.16fF $ **FLOATING
C1205 VDD.n272 VSS 0.01fF $ **FLOATING
C1206 VDD.n273 VSS 0.00fF $ **FLOATING
C1207 VDD.n274 VSS 0.00fF $ **FLOATING
C1208 VDD.n275 VSS 0.00fF $ **FLOATING
C1209 VDD.n276 VSS 0.00fF $ **FLOATING
C1210 VDD.n277 VSS 0.00fF $ **FLOATING
C1211 VDD.n278 VSS 0.00fF $ **FLOATING
C1212 VDD.n279 VSS 0.00fF $ **FLOATING
C1213 VDD.n280 VSS 0.00fF $ **FLOATING
C1214 VDD.n281 VSS 0.01fF $ **FLOATING
C1215 VDD.n282 VSS 0.00fF $ **FLOATING
C1216 VDD.n283 VSS 0.00fF $ **FLOATING
C1217 VDD.n284 VSS 0.00fF $ **FLOATING
C1218 VDD.n285 VSS 0.00fF $ **FLOATING
C1219 VDD.n286 VSS 0.00fF $ **FLOATING
C1220 VDD.n287 VSS 0.00fF $ **FLOATING
C1221 VDD.n288 VSS 0.00fF $ **FLOATING
C1222 VDD.n289 VSS 0.00fF $ **FLOATING
C1223 VDD.n290 VSS 0.00fF $ **FLOATING
C1224 VDD.n291 VSS 0.00fF $ **FLOATING
C1225 VDD.n292 VSS 0.00fF $ **FLOATING
C1226 VDD.n293 VSS 0.00fF $ **FLOATING
C1227 VDD.n294 VSS 0.00fF $ **FLOATING
C1228 VDD.n295 VSS 0.00fF $ **FLOATING
C1229 VDD.n296 VSS 0.00fF $ **FLOATING
C1230 VDD.n297 VSS 0.00fF $ **FLOATING
C1231 VDD.n298 VSS 0.00fF $ **FLOATING
C1232 VDD.n299 VSS 0.00fF $ **FLOATING
C1233 VDD.n300 VSS 0.00fF $ **FLOATING
C1234 VDD.n301 VSS 0.00fF $ **FLOATING
C1235 VDD.n302 VSS 0.00fF $ **FLOATING
C1236 VDD.n303 VSS 0.00fF $ **FLOATING
C1237 VDD.n304 VSS 0.00fF $ **FLOATING
C1238 VDD.n305 VSS 0.00fF $ **FLOATING
C1239 VDD.n306 VSS 0.00fF $ **FLOATING
C1240 VDD.n307 VSS 0.00fF $ **FLOATING
C1241 VDD.n308 VSS 0.00fF $ **FLOATING
C1242 VDD.n309 VSS 0.00fF $ **FLOATING
C1243 VDD.n310 VSS 0.00fF $ **FLOATING
C1244 VDD.n311 VSS 0.00fF $ **FLOATING
C1245 VDD.n312 VSS 0.00fF $ **FLOATING
C1246 VDD.n313 VSS 0.00fF $ **FLOATING
C1247 VDD.n314 VSS 0.00fF $ **FLOATING
C1248 VDD.n315 VSS 0.00fF $ **FLOATING
C1249 VDD.n316 VSS 0.00fF $ **FLOATING
C1250 VDD.n317 VSS 0.00fF $ **FLOATING
C1251 VDD.n318 VSS 0.00fF $ **FLOATING
C1252 VDD.n319 VSS 0.00fF $ **FLOATING
C1253 VDD.n320 VSS 0.00fF $ **FLOATING
C1254 VDD.n321 VSS 0.00fF $ **FLOATING
C1255 VDD.n322 VSS 0.00fF $ **FLOATING
C1256 VDD.n323 VSS 0.00fF $ **FLOATING
C1257 VDD.n324 VSS 0.00fF $ **FLOATING
C1258 VDD.n325 VSS 0.00fF $ **FLOATING
C1259 VDD.n326 VSS 0.00fF $ **FLOATING
C1260 VDD.n327 VSS 0.01fF $ **FLOATING
C1261 VDD.n328 VSS 0.00fF $ **FLOATING
C1262 VDD.n329 VSS 0.00fF $ **FLOATING
C1263 VDD.n330 VSS 0.00fF $ **FLOATING
C1264 VDD.n331 VSS 0.00fF $ **FLOATING
C1265 VDD.n332 VSS 0.00fF $ **FLOATING
C1266 VDD.n333 VSS 0.00fF $ **FLOATING
C1267 VDD.n334 VSS 0.00fF $ **FLOATING
C1268 VDD.n335 VSS 0.00fF $ **FLOATING
C1269 VDD.n336 VSS 0.00fF $ **FLOATING
C1270 VDD.n337 VSS 0.00fF $ **FLOATING
C1271 VDD.n338 VSS 0.01fF $ **FLOATING
C1272 VDD.n339 VSS 0.00fF $ **FLOATING
C1273 VDD.n340 VSS 0.00fF $ **FLOATING
C1274 VDD.n341 VSS 0.00fF $ **FLOATING
C1275 VDD.n342 VSS 0.00fF $ **FLOATING
C1276 VDD.n343 VSS 0.00fF $ **FLOATING
C1277 VDD.n344 VSS 0.00fF $ **FLOATING
C1278 VDD.n345 VSS 0.00fF $ **FLOATING
C1279 VDD.n346 VSS 0.00fF $ **FLOATING
C1280 VDD.n347 VSS 0.00fF $ **FLOATING
C1281 VDD.n348 VSS 0.00fF $ **FLOATING
C1282 VDD.n349 VSS 0.01fF $ **FLOATING
C1283 VDD.n350 VSS 0.00fF $ **FLOATING
C1284 VDD.n351 VSS 0.00fF $ **FLOATING
C1285 VDD.n352 VSS 0.00fF $ **FLOATING
C1286 VDD.n353 VSS 0.00fF $ **FLOATING
C1287 VDD.n354 VSS 0.00fF $ **FLOATING
C1288 VDD.n355 VSS 0.00fF $ **FLOATING
C1289 VDD.n356 VSS 0.00fF $ **FLOATING
C1290 VDD.n357 VSS 0.00fF $ **FLOATING
C1291 VDD.n358 VSS 0.00fF $ **FLOATING
C1292 VDD.n359 VSS 0.00fF $ **FLOATING
C1293 VDD.n360 VSS 0.00fF $ **FLOATING
C1294 VDD.n361 VSS 0.00fF $ **FLOATING
C1295 VDD.n362 VSS 0.00fF $ **FLOATING
C1296 VDD.n363 VSS 0.00fF $ **FLOATING
C1297 VDD.n364 VSS 0.00fF $ **FLOATING
C1298 VDD.n365 VSS 0.01fF $ **FLOATING
C1299 VDD.n366 VSS 0.01fF $ **FLOATING
C1300 VDD.n367 VSS 0.00fF $ **FLOATING
C1301 VDD.n368 VSS 0.00fF $ **FLOATING
C1302 VDD.n369 VSS 0.00fF $ **FLOATING
C1303 VDD.n370 VSS 0.00fF $ **FLOATING
C1304 VDD.n371 VSS 0.00fF $ **FLOATING
C1305 VDD.n372 VSS 0.00fF $ **FLOATING
C1306 VDD.n373 VSS 0.00fF $ **FLOATING
C1307 VDD.n374 VSS 0.00fF $ **FLOATING
C1308 VDD.n375 VSS 0.00fF $ **FLOATING
C1309 VDD.n376 VSS 0.00fF $ **FLOATING
C1310 VDD.n377 VSS 0.01fF $ **FLOATING
C1311 VDD.n378 VSS 0.00fF $ **FLOATING
C1312 VDD.n379 VSS 0.00fF $ **FLOATING
C1313 VDD.n380 VSS 0.00fF $ **FLOATING
C1314 VDD.n381 VSS 0.00fF $ **FLOATING
C1315 VDD.n382 VSS 0.00fF $ **FLOATING
C1316 VDD.n383 VSS 0.00fF $ **FLOATING
C1317 VDD.n384 VSS 0.00fF $ **FLOATING
C1318 VDD.n385 VSS 0.00fF $ **FLOATING
C1319 VDD.n386 VSS 0.00fF $ **FLOATING
C1320 VDD.n387 VSS 0.00fF $ **FLOATING
C1321 VDD.n388 VSS 0.01fF $ **FLOATING
C1322 VDD.n389 VSS 0.00fF $ **FLOATING
C1323 VDD.n390 VSS 0.00fF $ **FLOATING
C1324 VDD.n391 VSS 0.00fF $ **FLOATING
C1325 VDD.n392 VSS 0.00fF $ **FLOATING
C1326 VDD.n393 VSS 0.00fF $ **FLOATING
C1327 VDD.n394 VSS 0.00fF $ **FLOATING
C1328 VDD.n395 VSS 0.00fF $ **FLOATING
C1329 VDD.n396 VSS 0.00fF $ **FLOATING
C1330 VDD.n397 VSS 0.00fF $ **FLOATING
C1331 VDD.n398 VSS 0.00fF $ **FLOATING
C1332 VDD.n399 VSS 0.00fF $ **FLOATING
C1333 VDD.n400 VSS 0.00fF $ **FLOATING
C1334 VDD.n401 VSS 0.00fF $ **FLOATING
C1335 VDD.n402 VSS 0.00fF $ **FLOATING
C1336 VDD.n403 VSS 0.00fF $ **FLOATING
C1337 VDD.n404 VSS 0.00fF $ **FLOATING
C1338 VDD.n405 VSS 0.00fF $ **FLOATING
C1339 VDD.n406 VSS 0.00fF $ **FLOATING
C1340 VDD.n407 VSS 0.00fF $ **FLOATING
C1341 VDD.n408 VSS 0.00fF $ **FLOATING
C1342 VDD.n409 VSS 0.00fF $ **FLOATING
C1343 VDD.n410 VSS 0.00fF $ **FLOATING
C1344 VDD.n411 VSS 0.00fF $ **FLOATING
C1345 VDD.n412 VSS 0.00fF $ **FLOATING
C1346 VDD.n413 VSS 0.00fF $ **FLOATING
C1347 VDD.n414 VSS 0.00fF $ **FLOATING
C1348 VDD.n415 VSS 0.00fF $ **FLOATING
C1349 VDD.n416 VSS 0.00fF $ **FLOATING
C1350 VDD.n417 VSS 0.00fF $ **FLOATING
C1351 VDD.n418 VSS 0.00fF $ **FLOATING
C1352 VDD.n419 VSS 0.00fF $ **FLOATING
C1353 VDD.n420 VSS 0.00fF $ **FLOATING
C1354 VDD.n421 VSS 0.00fF $ **FLOATING
C1355 VDD.n422 VSS 0.00fF $ **FLOATING
C1356 VDD.n423 VSS 0.00fF $ **FLOATING
C1357 VDD.n424 VSS 0.00fF $ **FLOATING
C1358 VDD.n425 VSS 0.00fF $ **FLOATING
C1359 VDD.n426 VSS 0.00fF $ **FLOATING
C1360 VDD.n427 VSS 0.00fF $ **FLOATING
C1361 VDD.n428 VSS 0.00fF $ **FLOATING
C1362 VDD.n429 VSS 0.00fF $ **FLOATING
C1363 VDD.n430 VSS 0.01fF $ **FLOATING
C1364 VDD.n431 VSS 0.00fF $ **FLOATING
C1365 VDD.n432 VSS 0.00fF $ **FLOATING
C1366 VDD.n433 VSS 0.00fF $ **FLOATING
C1367 VDD.n434 VSS 0.00fF $ **FLOATING
C1368 VDD.n435 VSS 0.00fF $ **FLOATING
C1369 VDD.n436 VSS 0.00fF $ **FLOATING
C1370 VDD.n437 VSS 0.00fF $ **FLOATING
C1371 VDD.n438 VSS 0.00fF $ **FLOATING
C1372 VDD.n439 VSS 0.01fF $ **FLOATING
C1373 VDD.n440 VSS 0.00fF $ **FLOATING
C1374 VDD.n441 VSS 0.01fF $ **FLOATING
C1375 VDD.n442 VSS 1.25fF $ **FLOATING
C1376 VDD.n443 VSS 8.10fF $ **FLOATING
C1377 VDD.n444 VSS 0.03fF $ **FLOATING
C1378 VDD.n445 VSS 0.01fF $ **FLOATING
C1379 VDD.n446 VSS 0.00fF $ **FLOATING
C1380 VDD.n447 VSS 0.01fF $ **FLOATING
C1381 VDD.n448 VSS 0.01fF $ **FLOATING
C1382 VDD.n451 VSS 0.07fF $ **FLOATING
C1383 VDD.n452 VSS 0.01fF $ **FLOATING
C1384 VDD.n453 VSS 0.06fF $ **FLOATING
C1385 VDD.n454 VSS 0.64fF $ **FLOATING
C1386 VDD.n455 VSS 8.92fF $ **FLOATING
C1387 VDD.n456 VSS 0.86fF $ **FLOATING
C1388 VDD.n457 VSS 0.06fF $ **FLOATING
C1389 VDD.n458 VSS 0.14fF $ **FLOATING
C1390 VDD.n459 VSS 0.06fF $ **FLOATING
C1391 VDD.n460 VSS 0.13fF $ **FLOATING
C1392 VDD.n461 VSS 7.91fF $ **FLOATING
C1393 VDD.n462 VSS 0.07fF $ **FLOATING
C1394 VDD.n463 VSS 0.04fF $ **FLOATING
C1395 VDD.n464 VSS 0.13fF $ **FLOATING
C1396 VDD.n465 VSS 0.05fF $ **FLOATING
C1397 VDD.n466 VSS 0.13fF $ **FLOATING
C1398 VDD.n467 VSS 0.06fF $ **FLOATING
C1399 VDD.n468 VSS 0.13fF $ **FLOATING
C1400 VDD.n469 VSS 0.05fF $ **FLOATING
C1401 VDD.n470 VSS 0.13fF $ **FLOATING
C1402 VDD.n471 VSS 5.73fF $ **FLOATING
C1403 VDD.n472 VSS 0.07fF $ **FLOATING
C1404 VDD.n473 VSS 0.05fF $ **FLOATING
C1405 VDD.n474 VSS 0.13fF $ **FLOATING
C1406 VDD.n475 VSS 0.06fF $ **FLOATING
C1407 VDD.n476 VSS 0.13fF $ **FLOATING
C1408 VDD.n477 VSS 0.06fF $ **FLOATING
C1409 VDD.n478 VSS 0.13fF $ **FLOATING
C1410 VDD.n479 VSS 5.73fF $ **FLOATING
C1411 VDD.n480 VSS 0.06fF $ **FLOATING
C1412 VDD.n481 VSS 0.05fF $ **FLOATING
C1413 VDD.n482 VSS 0.13fF $ **FLOATING
C1414 VDD.n483 VSS 0.06fF $ **FLOATING
C1415 VDD.n484 VSS 0.13fF $ **FLOATING
C1416 VDD.n485 VSS 0.06fF $ **FLOATING
C1417 VDD.n486 VSS 0.13fF $ **FLOATING
C1418 VDD.n487 VSS 5.73fF $ **FLOATING
C1419 VDD.n488 VSS 0.06fF $ **FLOATING
C1420 VDD.n489 VSS 0.05fF $ **FLOATING
C1421 VDD.n490 VSS 0.13fF $ **FLOATING
C1422 VDD.n491 VSS 0.06fF $ **FLOATING
C1423 VDD.n492 VSS 0.13fF $ **FLOATING
C1424 VDD.n493 VSS 0.06fF $ **FLOATING
C1425 VDD.n494 VSS 0.13fF $ **FLOATING
C1426 VDD.n495 VSS 5.73fF $ **FLOATING
C1427 VDD.n496 VSS 0.07fF $ **FLOATING
C1428 VDD.n497 VSS 0.04fF $ **FLOATING
C1429 VDD.n498 VSS 0.13fF $ **FLOATING
C1430 VDD.n499 VSS 0.05fF $ **FLOATING
C1431 VDD.n500 VSS 0.13fF $ **FLOATING
C1432 VDD.n501 VSS 0.06fF $ **FLOATING
C1433 VDD.n502 VSS 0.13fF $ **FLOATING
C1434 VDD.n503 VSS 0.05fF $ **FLOATING
C1435 VDD.n504 VSS 0.13fF $ **FLOATING
C1436 VDD.n505 VSS 5.73fF $ **FLOATING
C1437 VDD.n506 VSS 0.07fF $ **FLOATING
C1438 VDD.n507 VSS 0.05fF $ **FLOATING
C1439 VDD.n508 VSS 0.13fF $ **FLOATING
C1440 VDD.n509 VSS 0.06fF $ **FLOATING
C1441 VDD.n510 VSS 0.13fF $ **FLOATING
C1442 VDD.n511 VSS 0.06fF $ **FLOATING
C1443 VDD.n512 VSS 0.13fF $ **FLOATING
C1444 VDD.n513 VSS 5.73fF $ **FLOATING
C1445 VDD.n514 VSS 0.06fF $ **FLOATING
C1446 VDD.n515 VSS 0.05fF $ **FLOATING
C1447 VDD.n516 VSS 0.13fF $ **FLOATING
C1448 VDD.n517 VSS 0.06fF $ **FLOATING
C1449 VDD.n518 VSS 0.13fF $ **FLOATING
C1450 VDD.n519 VSS 0.06fF $ **FLOATING
C1451 VDD.n520 VSS 0.13fF $ **FLOATING
C1452 VDD.n521 VSS 5.73fF $ **FLOATING
C1453 VDD.n522 VSS 0.06fF $ **FLOATING
C1454 VDD.n523 VSS 0.05fF $ **FLOATING
C1455 VDD.n524 VSS 0.13fF $ **FLOATING
C1456 VDD.n525 VSS 0.06fF $ **FLOATING
C1457 VDD.n526 VSS 0.13fF $ **FLOATING
C1458 VDD.n527 VSS 0.06fF $ **FLOATING
C1459 VDD.n528 VSS 0.13fF $ **FLOATING
C1460 VDD.n529 VSS 5.73fF $ **FLOATING
C1461 VDD.n530 VSS 0.07fF $ **FLOATING
C1462 VDD.n531 VSS 0.04fF $ **FLOATING
C1463 VDD.n532 VSS 0.13fF $ **FLOATING
C1464 VDD.n533 VSS 0.05fF $ **FLOATING
C1465 VDD.n534 VSS 0.13fF $ **FLOATING
C1466 VDD.n535 VSS 0.06fF $ **FLOATING
C1467 VDD.n536 VSS 0.13fF $ **FLOATING
C1468 VDD.n537 VSS 0.05fF $ **FLOATING
C1469 VDD.n538 VSS 0.13fF $ **FLOATING
C1470 VDD.n539 VSS 5.73fF $ **FLOATING
C1471 VDD.n540 VSS 0.07fF $ **FLOATING
C1472 VDD.n541 VSS 0.05fF $ **FLOATING
C1473 VDD.n542 VSS 0.13fF $ **FLOATING
C1474 VDD.n543 VSS 0.06fF $ **FLOATING
C1475 VDD.n544 VSS 0.13fF $ **FLOATING
C1476 VDD.n545 VSS 0.06fF $ **FLOATING
C1477 VDD.n546 VSS 0.13fF $ **FLOATING
C1478 VDD.n547 VSS 5.73fF $ **FLOATING
C1479 VDD.n548 VSS 0.06fF $ **FLOATING
C1480 VDD.n549 VSS 0.05fF $ **FLOATING
C1481 VDD.n550 VSS 0.13fF $ **FLOATING
C1482 VDD.n551 VSS 0.06fF $ **FLOATING
C1483 VDD.n552 VSS 0.13fF $ **FLOATING
C1484 VDD.n553 VSS 0.06fF $ **FLOATING
C1485 VDD.n554 VSS 0.13fF $ **FLOATING
C1486 VDD.n555 VSS 5.73fF $ **FLOATING
C1487 VDD.n556 VSS 0.06fF $ **FLOATING
C1488 VDD.n557 VSS 0.05fF $ **FLOATING
C1489 VDD.n558 VSS 0.13fF $ **FLOATING
C1490 VDD.n559 VSS 0.06fF $ **FLOATING
C1491 VDD.n560 VSS 0.13fF $ **FLOATING
C1492 VDD.n561 VSS 0.06fF $ **FLOATING
C1493 VDD.n562 VSS 0.13fF $ **FLOATING
C1494 VDD.n563 VSS 5.73fF $ **FLOATING
C1495 VDD.n564 VSS 0.07fF $ **FLOATING
C1496 VDD.n565 VSS 0.04fF $ **FLOATING
C1497 VDD.n566 VSS 0.13fF $ **FLOATING
C1498 VDD.n567 VSS 0.05fF $ **FLOATING
C1499 VDD.n568 VSS 0.13fF $ **FLOATING
C1500 VDD.n569 VSS 0.06fF $ **FLOATING
C1501 VDD.n570 VSS 0.13fF $ **FLOATING
C1502 VDD.n571 VSS 0.05fF $ **FLOATING
C1503 VDD.n572 VSS 0.13fF $ **FLOATING
C1504 VDD.n573 VSS 5.73fF $ **FLOATING
C1505 VDD.n574 VSS 0.07fF $ **FLOATING
C1506 VDD.n575 VSS 0.05fF $ **FLOATING
C1507 VDD.n576 VSS 0.13fF $ **FLOATING
C1508 VDD.n577 VSS 0.06fF $ **FLOATING
C1509 VDD.n578 VSS 0.13fF $ **FLOATING
C1510 VDD.n579 VSS 0.06fF $ **FLOATING
C1511 VDD.n580 VSS 0.13fF $ **FLOATING
C1512 VDD.n581 VSS 5.73fF $ **FLOATING
C1513 VDD.n582 VSS 0.06fF $ **FLOATING
C1514 VDD.n583 VSS 0.05fF $ **FLOATING
C1515 VDD.n584 VSS 0.13fF $ **FLOATING
C1516 VDD.n585 VSS 0.06fF $ **FLOATING
C1517 VDD.n586 VSS 0.13fF $ **FLOATING
C1518 VDD.n587 VSS 0.06fF $ **FLOATING
C1519 VDD.n588 VSS 0.11fF $ **FLOATING
C1520 VDD.n589 VSS 0.54fF $ **FLOATING
C1521 VDD.n590 VSS 5.73fF $ **FLOATING
C1522 VDD.n591 VSS 0.06fF $ **FLOATING
C1523 VDD.n592 VSS 0.05fF $ **FLOATING
C1524 VDD.n593 VSS 0.08fF $ **FLOATING
C1525 VDD.n594 VSS 0.06fF $ **FLOATING
C1526 VDD.n595 VSS 0.13fF $ **FLOATING
C1527 VDD.n596 VSS 0.06fF $ **FLOATING
C1528 VDD.n597 VSS 0.13fF $ **FLOATING
C1529 VDD.n598 VSS 5.73fF $ **FLOATING
C1530 VDD.n599 VSS 0.07fF $ **FLOATING
C1531 VDD.n600 VSS 0.04fF $ **FLOATING
C1532 VDD.n601 VSS 0.13fF $ **FLOATING
C1533 VDD.n602 VSS 0.05fF $ **FLOATING
C1534 VDD.n603 VSS 0.13fF $ **FLOATING
C1535 VDD.n604 VSS 0.06fF $ **FLOATING
C1536 VDD.n605 VSS 0.13fF $ **FLOATING
C1537 VDD.n606 VSS 0.05fF $ **FLOATING
C1538 VDD.n607 VSS 0.13fF $ **FLOATING
C1539 VDD.n608 VSS 5.73fF $ **FLOATING
C1540 VDD.n609 VSS 0.07fF $ **FLOATING
C1541 VDD.n610 VSS 0.05fF $ **FLOATING
C1542 VDD.n611 VSS 0.13fF $ **FLOATING
C1543 VDD.n612 VSS 0.06fF $ **FLOATING
C1544 VDD.n613 VSS 0.13fF $ **FLOATING
C1545 VDD.n614 VSS 0.06fF $ **FLOATING
C1546 VDD.n615 VSS 0.13fF $ **FLOATING
C1547 VDD.n616 VSS 7.60fF $ **FLOATING
C1548 VDD.n617 VSS 0.06fF $ **FLOATING
C1549 VDD.n618 VSS 0.05fF $ **FLOATING
C1550 VDD.n619 VSS 0.13fF $ **FLOATING
C1551 VDD.n620 VSS 0.06fF $ **FLOATING
C1552 VDD.n621 VSS 0.13fF $ **FLOATING
C1553 VDD.n622 VSS 0.36fF $ **FLOATING
C1554 VDD.n623 VSS 0.10fF $ **FLOATING
C1555 VDD.n624 VSS 0.26fF $ **FLOATING
C1556 VDD.n625 VSS 0.61fF $ **FLOATING
C1557 VDD.n626 VSS 0.06fF $ **FLOATING
C1558 VDD.n627 VSS 0.13fF $ **FLOATING
C1559 VDD.n628 VSS 0.13fF $ **FLOATING
C1560 VDD.n629 VSS 0.14fF $ **FLOATING
C1561 VDD.n630 VSS 0.05fF $ **FLOATING
C1562 VDD.n631 VSS 0.08fF $ **FLOATING
C1563 VDD.n632 VSS 1.02fF $ **FLOATING
C1564 VDD.t28 VSS 1.36fF
C1565 VDD.t22 VSS 2.02fF
C1566 VDD.t10 VSS 1.50fF
C1567 VDD.t1 VSS 2.02fF
C1568 VDD.t4 VSS 1.53fF
C1569 VDD.n633 VSS 1.02fF $ **FLOATING
C1570 VDD.n634 VSS 0.07fF $ **FLOATING
C1571 VDD.n635 VSS 0.05fF $ **FLOATING
C1572 VDD.n636 VSS 0.06fF $ **FLOATING
C1573 VDD.n637 VSS 0.13fF $ **FLOATING
C1574 VDD.n638 VSS 0.13fF $ **FLOATING
C1575 VDD.n639 VSS 0.13fF $ **FLOATING
C1576 VDD.n640 VSS 0.05fF $ **FLOATING
C1577 VDD.n641 VSS 0.06fF $ **FLOATING
C1578 VDD.n642 VSS 1.02fF $ **FLOATING
C1579 VDD.t13 VSS 1.69fF
C1580 VDD.t34 VSS 2.57fF
C1581 VDD.n643 VSS 0.14fF $ **FLOATING
C1582 VDD.n644 VSS 0.10fF $ **FLOATING
C1583 VDD.n645 VSS 0.07fF $ **FLOATING
C1584 VDD.n646 VSS 1.82fF $ **FLOATING
C1585 VDD.n647 VSS 0.38fF $ **FLOATING
C1586 VDD.n648 VSS 0.01fF $ **FLOATING
C1587 VDD.n649 VSS 0.00fF $ **FLOATING
C1588 VDD.n650 VSS 0.01fF $ **FLOATING
C1589 VDD.n651 VSS 0.01fF $ **FLOATING
C1590 VDD.n652 VSS 0.06fF $ **FLOATING
C1591 VDD.n653 VSS 0.01fF $ **FLOATING
C1592 VDD.n654 VSS 0.03fF $ **FLOATING
C1593 VDD.n655 VSS 0.01fF $ **FLOATING
C1594 VDD.n656 VSS 0.00fF $ **FLOATING
C1595 VDD.n657 VSS 0.01fF $ **FLOATING
C1596 VDD.n658 VSS 0.01fF $ **FLOATING
C1597 VDD.n659 VSS 0.09fF $ **FLOATING
C1598 VDD.n660 VSS 0.01fF $ **FLOATING
C1599 VDD.n661 VSS 0.07fF $ **FLOATING
C1600 VDD.n662 VSS 0.01fF $ **FLOATING
C1601 VDD.n663 VSS 0.07fF $ **FLOATING
C1602 VDD.n664 VSS 0.01fF $ **FLOATING
C1603 VDD.n665 VSS 0.07fF $ **FLOATING
C1604 VDD.n666 VSS 0.03fF $ **FLOATING
C1605 VDD.n667 VSS 0.13fF $ **FLOATING
C1606 VDD.n668 VSS 0.06fF $ **FLOATING
C1607 VDD.n669 VSS 5.73fF $ **FLOATING
C1608 VDD.n670 VSS 0.06fF $ **FLOATING
C1609 VDD.n671 VSS 0.13fF $ **FLOATING
C1610 VDD.n672 VSS 0.06fF $ **FLOATING
C1611 VDD.n673 VSS 0.13fF $ **FLOATING
C1612 VDD.n674 VSS 0.04fF $ **FLOATING
C1613 VDD.n675 VSS 5.73fF $ **FLOATING
C1614 VDD.n676 VSS 0.05fF $ **FLOATING
C1615 VDD.n677 VSS 0.06fF $ **FLOATING
C1616 VDD.n678 VSS 0.13fF $ **FLOATING
C1617 VDD.n679 VSS 0.06fF $ **FLOATING
C1618 VDD.n680 VSS 0.13fF $ **FLOATING
C1619 VDD.n681 VSS 0.07fF $ **FLOATING
C1620 VDD.n682 VSS 0.13fF $ **FLOATING
C1621 VDD.n683 VSS 0.07fF $ **FLOATING
C1622 VDD.n684 VSS 0.13fF $ **FLOATING
C1623 VDD.n685 VSS 0.06fF $ **FLOATING
C1624 VDD.n686 VSS 0.13fF $ **FLOATING
C1625 VDD.n687 VSS 0.05fF $ **FLOATING
C1626 VDD.n688 VSS 0.13fF $ **FLOATING
C1627 VDD.n689 VSS 0.06fF $ **FLOATING
C1628 VDD.n690 VSS 5.73fF $ **FLOATING
C1629 VDD.n691 VSS 0.05fF $ **FLOATING
C1630 VDD.n692 VSS 0.13fF $ **FLOATING
C1631 VDD.n693 VSS 0.06fF $ **FLOATING
C1632 VDD.n694 VSS 0.13fF $ **FLOATING
C1633 VDD.n695 VSS 0.05fF $ **FLOATING
C1634 VDD.n696 VSS 5.73fF $ **FLOATING
C1635 VDD.n697 VSS 0.06fF $ **FLOATING
C1636 VDD.n698 VSS 0.06fF $ **FLOATING
C1637 VDD.n699 VSS 0.13fF $ **FLOATING
C1638 VDD.n700 VSS 0.06fF $ **FLOATING
C1639 VDD.n701 VSS 0.13fF $ **FLOATING
C1640 VDD.n702 VSS 0.04fF $ **FLOATING
C1641 VDD.n703 VSS 5.73fF $ **FLOATING
C1642 VDD.n704 VSS 0.05fF $ **FLOATING
C1643 VDD.n705 VSS 0.06fF $ **FLOATING
C1644 VDD.n706 VSS 0.13fF $ **FLOATING
C1645 VDD.n707 VSS 0.06fF $ **FLOATING
C1646 VDD.n708 VSS 0.13fF $ **FLOATING
C1647 VDD.n709 VSS 0.07fF $ **FLOATING
C1648 VDD.n710 VSS 0.13fF $ **FLOATING
C1649 VDD.n711 VSS 0.07fF $ **FLOATING
C1650 VDD.n712 VSS 0.13fF $ **FLOATING
C1651 VDD.n713 VSS 5.73fF $ **FLOATING
C1652 VDD.n714 VSS 7.91fF $ **FLOATING
C1653 VDD.n715 VSS 8.92fF $ **FLOATING
C1654 VDD.n716 VSS 0.03fF $ **FLOATING
C1655 VDD.n717 VSS 0.01fF $ **FLOATING
C1656 VDD.n718 VSS 0.00fF $ **FLOATING
C1657 VDD.n719 VSS 0.01fF $ **FLOATING
C1658 VDD.n720 VSS 0.01fF $ **FLOATING
C1659 VDD.n723 VSS 0.07fF $ **FLOATING
C1660 VDD.n724 VSS 0.01fF $ **FLOATING
C1661 VDD.n725 VSS 0.06fF $ **FLOATING
C1662 VDD.n726 VSS 0.80fF $ **FLOATING
C1663 VDD.n727 VSS 0.75fF $ **FLOATING
C1664 VDD.n728 VSS 0.14fF $ **FLOATING
C1665 VDD.n729 VSS 0.06fF $ **FLOATING
C1666 VDD.n730 VSS 0.06fF $ **FLOATING
C1667 VDD.n731 VSS 0.04fF $ **FLOATING
C1668 VDD.n732 VSS 0.13fF $ **FLOATING
C1669 VDD.n733 VSS 0.13fF $ **FLOATING
C1670 VDD.n734 VSS 0.05fF $ **FLOATING
C1671 VDD.n735 VSS 0.06fF $ **FLOATING
C1672 VDD.n736 VSS 0.05fF $ **FLOATING
C1673 VDD.n737 VSS 0.13fF $ **FLOATING
C1674 VDD.n738 VSS 0.13fF $ **FLOATING
C1675 VDD.n739 VSS 0.05fF $ **FLOATING
C1676 VDD.n740 VSS 0.06fF $ **FLOATING
C1677 VDD.n741 VSS 0.06fF $ **FLOATING
C1678 VDD.n742 VSS 0.13fF $ **FLOATING
C1679 VDD.n743 VSS 0.13fF $ **FLOATING
C1680 VDD.n744 VSS 0.05fF $ **FLOATING
C1681 VDD.n745 VSS 0.06fF $ **FLOATING
C1682 VDD.n746 VSS 0.06fF $ **FLOATING
C1683 VDD.n747 VSS 0.13fF $ **FLOATING
C1684 VDD.n748 VSS 0.13fF $ **FLOATING
C1685 VDD.n749 VSS 0.13fF $ **FLOATING
C1686 VDD.n750 VSS 0.13fF $ **FLOATING
C1687 VDD.n751 VSS 0.06fF $ **FLOATING
C1688 VDD.n752 VSS 0.06fF $ **FLOATING
C1689 VDD.n753 VSS 5.73fF $ **FLOATING
C1690 VDD.n754 VSS 5.73fF $ **FLOATING
C1691 VDD.n755 VSS 0.07fF $ **FLOATING
C1692 VDD.n756 VSS 0.05fF $ **FLOATING
C1693 VDD.n757 VSS 0.13fF $ **FLOATING
C1694 VDD.n758 VSS 0.13fF $ **FLOATING
C1695 VDD.n759 VSS 0.13fF $ **FLOATING
C1696 VDD.n760 VSS 0.05fF $ **FLOATING
C1697 VDD.n761 VSS 0.07fF $ **FLOATING
C1698 VDD.n762 VSS 0.05fF $ **FLOATING
C1699 VDD.n763 VSS 0.06fF $ **FLOATING
C1700 VDD.n764 VSS 0.13fF $ **FLOATING
C1701 VDD.n765 VSS 0.13fF $ **FLOATING
C1702 VDD.n766 VSS 0.06fF $ **FLOATING
C1703 VDD.n767 VSS 0.13fF $ **FLOATING
C1704 VDD.n768 VSS 0.13fF $ **FLOATING
C1705 VDD.n769 VSS 0.13fF $ **FLOATING
C1706 VDD.n770 VSS 0.05fF $ **FLOATING
C1707 VDD.n771 VSS 0.06fF $ **FLOATING
C1708 VDD.n772 VSS 5.73fF $ **FLOATING
C1709 VDD.n773 VSS 5.73fF $ **FLOATING
C1710 VDD.n774 VSS 0.06fF $ **FLOATING
C1711 VDD.n775 VSS 0.06fF $ **FLOATING
C1712 VDD.n776 VSS 0.13fF $ **FLOATING
C1713 VDD.n777 VSS 0.13fF $ **FLOATING
C1714 VDD.n778 VSS 0.13fF $ **FLOATING
C1715 VDD.n779 VSS 0.04fF $ **FLOATING
C1716 VDD.n780 VSS 0.07fF $ **FLOATING
C1717 VDD.n781 VSS 0.05fF $ **FLOATING
C1718 VDD.n782 VSS 0.06fF $ **FLOATING
C1719 VDD.n783 VSS 0.13fF $ **FLOATING
C1720 VDD.n784 VSS 0.13fF $ **FLOATING
C1721 VDD.n785 VSS 0.13fF $ **FLOATING
C1722 VDD.n786 VSS 0.05fF $ **FLOATING
C1723 VDD.n787 VSS 0.07fF $ **FLOATING
C1724 VDD.n788 VSS 5.73fF $ **FLOATING
C1725 VDD.n789 VSS 5.73fF $ **FLOATING
C1726 VDD.n790 VSS 5.73fF $ **FLOATING
C1727 VDD.n791 VSS 5.73fF $ **FLOATING
C1728 VDD.n792 VSS 5.73fF $ **FLOATING
C1729 VDD.n793 VSS 0.06fF $ **FLOATING
C1730 VDD.n794 VSS 0.06fF $ **FLOATING
C1731 VDD.n795 VSS 0.13fF $ **FLOATING
C1732 VDD.n796 VSS 0.13fF $ **FLOATING
C1733 VDD.n797 VSS 0.13fF $ **FLOATING
C1734 VDD.n798 VSS 0.06fF $ **FLOATING
C1735 VDD.n799 VSS 0.06fF $ **FLOATING
C1736 VDD.n800 VSS 0.05fF $ **FLOATING
C1737 VDD.n801 VSS 0.13fF $ **FLOATING
C1738 VDD.n802 VSS 0.13fF $ **FLOATING
C1739 VDD.n803 VSS 0.06fF $ **FLOATING
C1740 VDD.n804 VSS 0.06fF $ **FLOATING
C1741 VDD.n805 VSS 0.04fF $ **FLOATING
C1742 VDD.n806 VSS 0.13fF $ **FLOATING
C1743 VDD.n807 VSS 0.13fF $ **FLOATING
C1744 VDD.n808 VSS 0.05fF $ **FLOATING
C1745 VDD.n809 VSS 0.06fF $ **FLOATING
C1746 VDD.n810 VSS 0.05fF $ **FLOATING
C1747 VDD.n811 VSS 0.13fF $ **FLOATING
C1748 VDD.n812 VSS 0.13fF $ **FLOATING
C1749 VDD.n813 VSS 0.05fF $ **FLOATING
C1750 VDD.n814 VSS 0.06fF $ **FLOATING
C1751 VDD.n815 VSS 0.06fF $ **FLOATING
C1752 VDD.n816 VSS 0.13fF $ **FLOATING
C1753 VDD.n817 VSS 0.13fF $ **FLOATING
C1754 VDD.n818 VSS 0.05fF $ **FLOATING
C1755 VDD.n819 VSS 0.06fF $ **FLOATING
C1756 VDD.n820 VSS 0.06fF $ **FLOATING
C1757 VDD.n821 VSS 0.13fF $ **FLOATING
C1758 VDD.n822 VSS 0.13fF $ **FLOATING
C1759 VDD.n823 VSS 0.13fF $ **FLOATING
C1760 VDD.n824 VSS 0.13fF $ **FLOATING
C1761 VDD.n825 VSS 0.06fF $ **FLOATING
C1762 VDD.n826 VSS 0.06fF $ **FLOATING
C1763 VDD.n827 VSS 5.73fF $ **FLOATING
C1764 VDD.n828 VSS 5.73fF $ **FLOATING
C1765 VDD.n829 VSS 0.07fF $ **FLOATING
C1766 VDD.n830 VSS 0.05fF $ **FLOATING
C1767 VDD.n831 VSS 0.10fF $ **FLOATING
C1768 VDD.n832 VSS 9.74fF $ **FLOATING
C1769 VDD.n833 VSS 0.10fF $ **FLOATING
C1770 VDD.n834 VSS 0.13fF $ **FLOATING
C1771 VDD.n835 VSS 0.05fF $ **FLOATING
C1772 VDD.n836 VSS 0.07fF $ **FLOATING
C1773 VDD.n837 VSS 0.05fF $ **FLOATING
C1774 VDD.n838 VSS 0.06fF $ **FLOATING
C1775 VDD.n839 VSS 0.13fF $ **FLOATING
C1776 VDD.n840 VSS 0.13fF $ **FLOATING
C1777 VDD.n841 VSS 0.13fF $ **FLOATING
C1778 VDD.n842 VSS 0.05fF $ **FLOATING
C1779 VDD.n843 VSS 0.06fF $ **FLOATING
C1780 VDD.n844 VSS 7.60fF $ **FLOATING
C1781 VDD.n845 VSS 0.36fF $ **FLOATING
C1782 VDD.n846 VSS 0.10fF $ **FLOATING
C1783 VDD.n847 VSS 1.85fF $ **FLOATING
C1784 VDD.n848 VSS 0.44fF $ **FLOATING
C1785 VDD.n849 VSS 0.01fF $ **FLOATING
C1786 VDD.n850 VSS 0.00fF $ **FLOATING
C1787 VDD.n851 VSS 0.01fF $ **FLOATING
C1788 VDD.n852 VSS 0.01fF $ **FLOATING
C1789 VDD.n853 VSS 0.06fF $ **FLOATING
C1790 VDD.n854 VSS 0.01fF $ **FLOATING
C1791 VDD.n855 VSS 0.03fF $ **FLOATING
C1792 VDD.n856 VSS 0.01fF $ **FLOATING
C1793 VDD.n857 VSS 0.00fF $ **FLOATING
C1794 VDD.n858 VSS 0.01fF $ **FLOATING
C1795 VDD.n859 VSS 0.01fF $ **FLOATING
C1796 VDD.n860 VSS 0.09fF $ **FLOATING
C1797 VDD.n861 VSS 0.01fF $ **FLOATING
C1798 VDD.n862 VSS 0.07fF $ **FLOATING
C1799 VDD.n863 VSS 0.01fF $ **FLOATING
C1800 VDD.n864 VSS 0.07fF $ **FLOATING
C1801 VDD.n865 VSS 0.01fF $ **FLOATING
C1802 VDD.n866 VSS 0.07fF $ **FLOATING
C1803 VDD.n867 VSS 0.03fF $ **FLOATING
C1804 VDD.n868 VSS 1.94fF $ **FLOATING
C1805 VDD.n869 VSS 0.06fF $ **FLOATING
C1806 VDD.n870 VSS 8.01fF $ **FLOATING
C1807 VDD.n871 VSS 0.06fF $ **FLOATING
C1808 VDD.n872 VSS 0.13fF $ **FLOATING
C1809 VDD.n873 VSS 0.06fF $ **FLOATING
C1810 VDD.n874 VSS 0.03fF $ **FLOATING
C1811 VDD.n875 VSS 0.01fF $ **FLOATING
C1812 VDD.n876 VSS 0.00fF $ **FLOATING
C1813 VDD.n877 VSS 0.01fF $ **FLOATING
C1814 VDD.n878 VSS 0.01fF $ **FLOATING
C1815 VDD.n881 VSS 0.07fF $ **FLOATING
C1816 VDD.n882 VSS 0.01fF $ **FLOATING
C1817 VDD.n883 VSS 0.06fF $ **FLOATING
C1818 VDD.n884 VSS 2.77fF $ **FLOATING
C1819 VDD.n885 VSS 0.57fF $ **FLOATING
C1820 VDD.n886 VSS 9.32fF $ **FLOATING
C1821 VDD.n887 VSS 0.05fF $ **FLOATING
C1822 VDD.n888 VSS 0.14fF $ **FLOATING
C1823 VDD.n889 VSS 0.13fF $ **FLOATING
C1824 VDD.n890 VSS 0.13fF $ **FLOATING
C1825 VDD.n891 VSS 0.05fF $ **FLOATING
C1826 VDD.n892 VSS 0.07fF $ **FLOATING
C1827 VDD.n893 VSS 0.05fF $ **FLOATING
C1828 VDD.n894 VSS 0.06fF $ **FLOATING
C1829 VDD.n895 VSS 0.13fF $ **FLOATING
C1830 VDD.n896 VSS 0.13fF $ **FLOATING
C1831 VDD.n897 VSS 0.08fF $ **FLOATING
C1832 VDD.n898 VSS 0.13fF $ **FLOATING
C1833 VDD.n899 VSS 0.05fF $ **FLOATING
C1834 VDD.n900 VSS 0.06fF $ **FLOATING
C1835 VDD.n901 VSS 7.60fF $ **FLOATING
C1836 VDD.n902 VSS 0.36fF $ **FLOATING
C1837 VDD.n903 VSS 0.10fF $ **FLOATING
C1838 VDD.n904 VSS 0.83fF $ **FLOATING
C1839 VDD.n905 VSS 0.44fF $ **FLOATING
C1840 VDD.n906 VSS 0.01fF $ **FLOATING
C1841 VDD.n907 VSS 0.00fF $ **FLOATING
C1842 VDD.n908 VSS 0.01fF $ **FLOATING
C1843 VDD.n909 VSS 0.01fF $ **FLOATING
C1844 VDD.n910 VSS 0.06fF $ **FLOATING
C1845 VDD.n911 VSS 0.01fF $ **FLOATING
C1846 VDD.n912 VSS 0.03fF $ **FLOATING
C1847 VDD.n913 VSS 0.01fF $ **FLOATING
C1848 VDD.n914 VSS 0.00fF $ **FLOATING
C1849 VDD.n915 VSS 0.01fF $ **FLOATING
C1850 VDD.n916 VSS 0.01fF $ **FLOATING
C1851 VDD.n917 VSS 0.09fF $ **FLOATING
C1852 VDD.n918 VSS 0.01fF $ **FLOATING
C1853 VDD.n919 VSS 0.07fF $ **FLOATING
C1854 VDD.n920 VSS 0.01fF $ **FLOATING
C1855 VDD.n922 VSS 0.07fF $ **FLOATING
C1856 VDD.n923 VSS 0.01fF $ **FLOATING
C1857 VDD.n924 VSS 0.07fF $ **FLOATING
C1858 VDD.n925 VSS 0.03fF $ **FLOATING
C1859 VDD.n926 VSS 0.03fF $ **FLOATING
C1860 VDD.n927 VSS 0.01fF $ **FLOATING
C1861 VDD.n928 VSS 0.00fF $ **FLOATING
C1862 VDD.n929 VSS 0.01fF $ **FLOATING
C1863 VDD.n930 VSS 0.01fF $ **FLOATING
C1864 VDD.n933 VSS 0.07fF $ **FLOATING
C1865 VDD.n934 VSS 0.01fF $ **FLOATING
C1866 VDD.n935 VSS 0.06fF $ **FLOATING
C1867 VDD.n936 VSS 2.77fF $ **FLOATING
C1868 VDD.n937 VSS 32.87fF $ **FLOATING
C1869 VDD.n938 VSS 26.20fF $ **FLOATING
C1870 VDD.n939 VSS 27.34fF $ **FLOATING
C1871 VDD.n940 VSS 1.86fF $ **FLOATING
C1872 VDD.n941 VSS 7.34fF $ **FLOATING
C1873 VDD.n942 VSS 1.66fF $ **FLOATING
C1874 VDD.n943 VSS 0.01fF $ **FLOATING
C1875 VDD.n944 VSS 0.00fF $ **FLOATING
C1876 VDD.n945 VSS 0.01fF $ **FLOATING
C1877 VDD.n946 VSS 0.01fF $ **FLOATING
C1878 VDD.n947 VSS 0.06fF $ **FLOATING
C1879 VDD.n948 VSS 0.01fF $ **FLOATING
C1880 VDD.n949 VSS 0.03fF $ **FLOATING
C1881 VDD.n950 VSS 0.01fF $ **FLOATING
C1882 VDD.n951 VSS 0.00fF $ **FLOATING
C1883 VDD.n952 VSS 0.01fF $ **FLOATING
C1884 VDD.n953 VSS 0.01fF $ **FLOATING
C1885 VDD.n954 VSS 0.09fF $ **FLOATING
C1886 VDD.n955 VSS 0.01fF $ **FLOATING
C1887 VDD.n956 VSS 0.07fF $ **FLOATING
C1888 VDD.n957 VSS 0.01fF $ **FLOATING
C1889 VDD.n959 VSS 0.07fF $ **FLOATING
C1890 VDD.n960 VSS 0.01fF $ **FLOATING
C1891 VDD.n961 VSS 0.07fF $ **FLOATING
C1892 VDD.n962 VSS 0.03fF $ **FLOATING
C1893 VDD.n963 VSS 0.03fF $ **FLOATING
C1894 VDD.n964 VSS 0.01fF $ **FLOATING
C1895 VDD.n965 VSS 0.00fF $ **FLOATING
C1896 VDD.n966 VSS 0.01fF $ **FLOATING
C1897 VDD.n967 VSS 0.01fF $ **FLOATING
C1898 VDD.n970 VSS 0.07fF $ **FLOATING
C1899 VDD.n971 VSS 0.01fF $ **FLOATING
C1900 VDD.n972 VSS 0.06fF $ **FLOATING
C1901 VDD.n973 VSS 2.77fF $ **FLOATING
C1902 VDD.n974 VSS 2.40fF $ **FLOATING
C1903 VDD.n975 VSS 0.01fF $ **FLOATING
C1904 VDD.n976 VSS 0.00fF $ **FLOATING
C1905 VDD.n977 VSS 0.01fF $ **FLOATING
C1906 VDD.n978 VSS 0.01fF $ **FLOATING
C1907 VDD.n979 VSS 0.06fF $ **FLOATING
C1908 VDD.n980 VSS 0.01fF $ **FLOATING
C1909 VDD.n981 VSS 0.03fF $ **FLOATING
C1910 VDD.n982 VSS 0.01fF $ **FLOATING
C1911 VDD.n983 VSS 0.00fF $ **FLOATING
C1912 VDD.n984 VSS 0.01fF $ **FLOATING
C1913 VDD.n985 VSS 0.01fF $ **FLOATING
C1914 VDD.n986 VSS 0.09fF $ **FLOATING
C1915 VDD.n987 VSS 0.01fF $ **FLOATING
C1916 VDD.n988 VSS 0.07fF $ **FLOATING
C1917 VDD.n989 VSS 0.01fF $ **FLOATING
C1918 VDD.n990 VSS 0.07fF $ **FLOATING
C1919 VDD.n991 VSS 0.01fF $ **FLOATING
C1920 VDD.n992 VSS 0.07fF $ **FLOATING
C1921 VDD.n993 VSS 0.03fF $ **FLOATING
C1922 VDD.n994 VSS 0.03fF $ **FLOATING
C1923 VDD.n995 VSS 0.01fF $ **FLOATING
C1924 VDD.n996 VSS 0.00fF $ **FLOATING
C1925 VDD.n997 VSS 0.01fF $ **FLOATING
C1926 VDD.n998 VSS 0.01fF $ **FLOATING
C1927 VDD.n1001 VSS 0.07fF $ **FLOATING
C1928 VDD.n1002 VSS 0.01fF $ **FLOATING
C1929 VDD.n1003 VSS 0.06fF $ **FLOATING
C1930 VDD.n1004 VSS 2.77fF $ **FLOATING
C1931 VDD.n1005 VSS 2.84fF $ **FLOATING
C1932 VDD.n1006 VSS 0.01fF $ **FLOATING
C1933 VDD.n1007 VSS 0.00fF $ **FLOATING
C1934 VDD.n1008 VSS 0.01fF $ **FLOATING
C1935 VDD.n1009 VSS 0.01fF $ **FLOATING
C1936 VDD.n1010 VSS 0.06fF $ **FLOATING
C1937 VDD.n1011 VSS 0.01fF $ **FLOATING
C1938 VDD.n1012 VSS 0.03fF $ **FLOATING
C1939 VDD.n1013 VSS 0.01fF $ **FLOATING
C1940 VDD.n1014 VSS 0.00fF $ **FLOATING
C1941 VDD.n1015 VSS 0.01fF $ **FLOATING
C1942 VDD.n1016 VSS 0.01fF $ **FLOATING
C1943 VDD.n1017 VSS 0.09fF $ **FLOATING
C1944 VDD.n1018 VSS 0.01fF $ **FLOATING
C1945 VDD.n1019 VSS 0.07fF $ **FLOATING
C1946 VDD.n1020 VSS 0.01fF $ **FLOATING
C1947 VDD.n1022 VSS 0.07fF $ **FLOATING
C1948 VDD.n1023 VSS 0.01fF $ **FLOATING
C1949 VDD.n1024 VSS 0.07fF $ **FLOATING
C1950 VDD.n1025 VSS 0.03fF $ **FLOATING
C1951 VDD.n1026 VSS 0.03fF $ **FLOATING
C1952 VDD.n1027 VSS 0.01fF $ **FLOATING
C1953 VDD.n1028 VSS 0.00fF $ **FLOATING
C1954 VDD.n1029 VSS 0.01fF $ **FLOATING
C1955 VDD.n1030 VSS 0.01fF $ **FLOATING
C1956 VDD.n1033 VSS 0.07fF $ **FLOATING
C1957 VDD.n1034 VSS 0.01fF $ **FLOATING
C1958 VDD.n1035 VSS 0.06fF $ **FLOATING
C1959 VDD.n1036 VSS 0.80fF $ **FLOATING
C1960 VDD.n1037 VSS 3.28fF $ **FLOATING
C1961 VDD.n1038 VSS 0.01fF $ **FLOATING
C1962 VDD.n1039 VSS 0.00fF $ **FLOATING
C1963 VDD.n1040 VSS 0.01fF $ **FLOATING
C1964 VDD.n1041 VSS 0.01fF $ **FLOATING
C1965 VDD.n1042 VSS 0.06fF $ **FLOATING
C1966 VDD.n1043 VSS 0.01fF $ **FLOATING
C1967 VDD.n1044 VSS 0.03fF $ **FLOATING
C1968 VDD.n1045 VSS 0.01fF $ **FLOATING
C1969 VDD.n1046 VSS 0.00fF $ **FLOATING
C1970 VDD.n1047 VSS 0.01fF $ **FLOATING
C1971 VDD.n1048 VSS 0.01fF $ **FLOATING
C1972 VDD.n1049 VSS 0.09fF $ **FLOATING
C1973 VDD.n1050 VSS 0.01fF $ **FLOATING
C1974 VDD.n1051 VSS 0.07fF $ **FLOATING
C1975 VDD.n1052 VSS 0.01fF $ **FLOATING
C1976 VDD.n1053 VSS 0.07fF $ **FLOATING
C1977 VDD.n1054 VSS 0.01fF $ **FLOATING
C1978 VDD.n1055 VSS 0.07fF $ **FLOATING
C1979 VDD.n1056 VSS 0.03fF $ **FLOATING
C1980 VDD.n1057 VSS 0.03fF $ **FLOATING
C1981 VDD.n1058 VSS 0.01fF $ **FLOATING
C1982 VDD.n1059 VSS 0.00fF $ **FLOATING
C1983 VDD.n1060 VSS 0.01fF $ **FLOATING
C1984 VDD.n1061 VSS 0.01fF $ **FLOATING
C1985 VDD.n1064 VSS 0.07fF $ **FLOATING
C1986 VDD.n1065 VSS 0.01fF $ **FLOATING
C1987 VDD.n1066 VSS 0.06fF $ **FLOATING
C1988 VDD.n1067 VSS 1.05fF $ **FLOATING
C1989 VDD.n1068 VSS 3.81fF $ **FLOATING
C1990 VDD.n1069 VSS 0.01fF $ **FLOATING
C1991 VDD.n1070 VSS 0.00fF $ **FLOATING
C1992 VDD.n1071 VSS 0.01fF $ **FLOATING
C1993 VDD.n1072 VSS 0.01fF $ **FLOATING
C1994 VDD.n1073 VSS 0.06fF $ **FLOATING
C1995 VDD.n1074 VSS 0.01fF $ **FLOATING
C1996 VDD.n1075 VSS 3.99fF $ **FLOATING
C1997 VDD.n1076 VSS 3.99fF $ **FLOATING
C1998 VDD.n1077 VSS 0.07fF $ **FLOATING
C1999 VDD.n1078 VSS 0.01fF $ **FLOATING
C2000 VDD.n1080 VSS 0.07fF $ **FLOATING
C2001 VDD.n1081 VSS 0.01fF $ **FLOATING
C2002 VDD.n1082 VSS 0.07fF $ **FLOATING
C2003 VDD.n1083 VSS 0.01fF $ **FLOATING
C2004 VDD.n1084 VSS 0.06fF $ **FLOATING
C2005 VDD.n1086 VSS 3.99fF $ **FLOATING
C2006 VDD.n1087 VSS 3.99fF $ **FLOATING
C2007 VDD.n1088 VSS 0.07fF $ **FLOATING
C2008 VDD.n1089 VSS 0.01fF $ **FLOATING
C2009 VDD.n1090 VSS 0.07fF $ **FLOATING
C2010 VDD.n1091 VSS 0.01fF $ **FLOATING
C2011 VDD.n1092 VSS 0.07fF $ **FLOATING
C2012 VDD.n1093 VSS 0.01fF $ **FLOATING
C2013 VDD.n1094 VSS 0.06fF $ **FLOATING
C2014 VDD.n1096 VSS 3.99fF $ **FLOATING
C2015 VDD.n1097 VSS 3.99fF $ **FLOATING
C2016 VDD.n1098 VSS 0.07fF $ **FLOATING
C2017 VDD.n1099 VSS 0.01fF $ **FLOATING
C2018 VDD.n1101 VSS 0.07fF $ **FLOATING
C2019 VDD.n1102 VSS 0.01fF $ **FLOATING
C2020 VDD.n1103 VSS 0.07fF $ **FLOATING
C2021 VDD.n1104 VSS 0.01fF $ **FLOATING
C2022 VDD.n1105 VSS 0.06fF $ **FLOATING
C2023 VDD.n1107 VSS 3.99fF $ **FLOATING
C2024 VDD.n1108 VSS 3.99fF $ **FLOATING
C2025 VDD.n1109 VSS 0.07fF $ **FLOATING
C2026 VDD.n1110 VSS 0.01fF $ **FLOATING
C2027 VDD.n1111 VSS 0.07fF $ **FLOATING
C2028 VDD.n1112 VSS 0.01fF $ **FLOATING
C2029 VDD.n1113 VSS 0.07fF $ **FLOATING
C2030 VDD.n1114 VSS 0.01fF $ **FLOATING
C2031 VDD.n1115 VSS 0.06fF $ **FLOATING
C2032 VDD.n1117 VSS 3.99fF $ **FLOATING
C2033 VDD.n1118 VSS 3.99fF $ **FLOATING
C2034 VDD.n1119 VSS 0.07fF $ **FLOATING
C2035 VDD.n1120 VSS 0.01fF $ **FLOATING
C2036 VDD.n1121 VSS 0.07fF $ **FLOATING
C2037 VDD.n1122 VSS 0.01fF $ **FLOATING
C2038 VDD.n1123 VSS 0.07fF $ **FLOATING
C2039 VDD.n1124 VSS 0.01fF $ **FLOATING
C2040 VDD.n1125 VSS 0.06fF $ **FLOATING
C2041 VDD.n1127 VSS 3.99fF $ **FLOATING
C2042 VDD.n1128 VSS 3.99fF $ **FLOATING
C2043 VDD.n1129 VSS 0.07fF $ **FLOATING
C2044 VDD.n1130 VSS 0.01fF $ **FLOATING
C2045 VDD.n1132 VSS 0.07fF $ **FLOATING
C2046 VDD.n1133 VSS 0.01fF $ **FLOATING
C2047 VDD.n1134 VSS 0.07fF $ **FLOATING
C2048 VDD.n1135 VSS 0.01fF $ **FLOATING
C2049 VDD.n1136 VSS 0.06fF $ **FLOATING
C2050 VDD.n1138 VSS 3.99fF $ **FLOATING
C2051 VDD.n1139 VSS 3.99fF $ **FLOATING
C2052 VDD.n1140 VSS 0.07fF $ **FLOATING
C2053 VDD.n1141 VSS 0.01fF $ **FLOATING
C2054 VDD.n1143 VSS 0.07fF $ **FLOATING
C2055 VDD.n1144 VSS 0.01fF $ **FLOATING
C2056 VDD.n1145 VSS 0.07fF $ **FLOATING
C2057 VDD.n1146 VSS 0.01fF $ **FLOATING
C2058 VDD.n1147 VSS 0.06fF $ **FLOATING
C2059 VDD.n1149 VSS 3.99fF $ **FLOATING
C2060 VDD.n1150 VSS 3.99fF $ **FLOATING
C2061 VDD.n1151 VSS 0.07fF $ **FLOATING
C2062 VDD.n1152 VSS 0.01fF $ **FLOATING
C2063 VDD.n1154 VSS 0.07fF $ **FLOATING
C2064 VDD.n1155 VSS 0.01fF $ **FLOATING
C2065 VDD.n1156 VSS 0.07fF $ **FLOATING
C2066 VDD.n1157 VSS 0.01fF $ **FLOATING
C2067 VDD.n1158 VSS 0.06fF $ **FLOATING
C2068 VDD.n1160 VSS 3.99fF $ **FLOATING
C2069 VDD.n1161 VSS 3.99fF $ **FLOATING
C2070 VDD.n1162 VSS 0.07fF $ **FLOATING
C2071 VDD.n1163 VSS 0.01fF $ **FLOATING
C2072 VDD.n1165 VSS 0.07fF $ **FLOATING
C2073 VDD.n1166 VSS 0.01fF $ **FLOATING
C2074 VDD.n1167 VSS 0.07fF $ **FLOATING
C2075 VDD.n1168 VSS 0.01fF $ **FLOATING
C2076 VDD.n1169 VSS 0.06fF $ **FLOATING
C2077 VDD.n1170 VSS 0.01fF $ **FLOATING
C2078 VDD.n1171 VSS 0.01fF $ **FLOATING
C2079 VDD.n1172 VSS 0.00fF $ **FLOATING
C2080 VDD.n1173 VSS 0.01fF $ **FLOATING
C2081 VDD.n1174 VSS 0.01fF $ **FLOATING
C2082 VDD.n1175 VSS 0.06fF $ **FLOATING
C2083 VDD.n1176 VSS 0.03fF $ **FLOATING
C2084 VDD.n1177 VSS 0.44fF $ **FLOATING
C2085 VDD.n1178 VSS 0.26fF $ **FLOATING
C2086 VDD.n1179 VSS 0.10fF $ **FLOATING
C2087 VDD.n1180 VSS 0.06fF $ **FLOATING
C2088 VDD.n1181 VSS 0.05fF $ **FLOATING
C2089 VDD.n1182 VSS 0.10fF $ **FLOATING
C2090 VDD.n1183 VSS 1.32fF $ **FLOATING
C2091 VDD.n1184 VSS 0.48fF $ **FLOATING
C2092 VDD.n1185 VSS 0.84fF $ **FLOATING
C2093 VDD.n1186 VSS 0.10fF $ **FLOATING
C2094 VDD.n1187 VSS 0.06fF $ **FLOATING
C2095 VDD.n1188 VSS 0.05fF $ **FLOATING
C2096 VDD.n1189 VSS 0.13fF $ **FLOATING
C2097 VDD.n1190 VSS 0.09fF $ **FLOATING
C2098 VDD.n1191 VSS 1.37fF $ **FLOATING
C2099 VDD.n1192 VSS 0.40fF $ **FLOATING
C2100 VDD.n1193 VSS 0.80fF $ **FLOATING
C2101 VDD.n1194 VSS 0.01fF $ **FLOATING
C2102 VDD.n1195 VSS 0.00fF $ **FLOATING
C2103 VDD.n1196 VSS 0.01fF $ **FLOATING
C2104 VDD.n1197 VSS 0.01fF $ **FLOATING
C2105 VDD.n1198 VSS 0.06fF $ **FLOATING
C2106 VDD.n1199 VSS 0.01fF $ **FLOATING
C2107 VDD.n1200 VSS 0.07fF $ **FLOATING
C2108 VDD.n1201 VSS 0.01fF $ **FLOATING
C2109 VDD.n1202 VSS 0.07fF $ **FLOATING
C2110 VDD.n1203 VSS 0.01fF $ **FLOATING
C2111 VDD.n1204 VSS 0.04fF $ **FLOATING
C2112 VDD.n1205 VSS 0.01fF $ **FLOATING
C2113 VDD.n1206 VSS 0.04fF $ **FLOATING
C2114 VDD.n1207 VSS 0.00fF $ **FLOATING
C2115 VDD.n1208 VSS 0.06fF $ **FLOATING
C2116 VDD.n1210 VSS 3.99fF $ **FLOATING
C2117 VDD.n1211 VSS 3.99fF $ **FLOATING
C2118 VDD.n1213 VSS 0.06fF $ **FLOATING
C2119 VDD.n1215 VSS 3.99fF $ **FLOATING
C2120 VDD.n1216 VSS 3.99fF $ **FLOATING
C2121 VDD.n1218 VSS 0.06fF $ **FLOATING
C2122 VDD.n1220 VSS 3.99fF $ **FLOATING
C2123 VDD.n1221 VSS 3.99fF $ **FLOATING
C2124 VDD.n1223 VSS 0.06fF $ **FLOATING
C2125 VDD.n1225 VSS 3.99fF $ **FLOATING
C2126 VDD.n1226 VSS 3.99fF $ **FLOATING
C2127 VDD.n1228 VSS 0.06fF $ **FLOATING
C2128 VDD.n1230 VSS 3.99fF $ **FLOATING
C2129 VDD.n1231 VSS 3.99fF $ **FLOATING
C2130 VDD.n1233 VSS 0.06fF $ **FLOATING
C2131 VDD.n1235 VSS 3.99fF $ **FLOATING
C2132 VDD.n1236 VSS 3.99fF $ **FLOATING
C2133 VDD.n1238 VSS 0.06fF $ **FLOATING
C2134 VDD.n1240 VSS 3.99fF $ **FLOATING
C2135 VDD.n1241 VSS 3.99fF $ **FLOATING
C2136 VDD.n1243 VSS 0.06fF $ **FLOATING
C2137 VDD.n1245 VSS 3.99fF $ **FLOATING
C2138 VDD.n1246 VSS 3.99fF $ **FLOATING
C2139 VDD.n1248 VSS 0.06fF $ **FLOATING
C2140 VDD.n1250 VSS 3.99fF $ **FLOATING
C2141 VDD.n1251 VSS 3.99fF $ **FLOATING
C2142 VDD.n1253 VSS 0.07fF $ **FLOATING
C2143 VDD.n1254 VSS 0.01fF $ **FLOATING
C2144 VDD.n1255 VSS 0.03fF $ **FLOATING
C2145 VDD.n1256 VSS 0.04fF $ **FLOATING
C2146 VDD.n1257 VSS 0.01fF $ **FLOATING
C2147 VDD.n1258 VSS 0.07fF $ **FLOATING
C2148 VDD.n1259 VSS 0.01fF $ **FLOATING
C2149 VDD.n1260 VSS 0.03fF $ **FLOATING
C2150 VDD.n1261 VSS 0.04fF $ **FLOATING
C2151 VDD.n1262 VSS 0.01fF $ **FLOATING
C2152 VDD.n1263 VSS 0.07fF $ **FLOATING
C2153 VDD.n1264 VSS 0.01fF $ **FLOATING
C2154 VDD.n1265 VSS 0.03fF $ **FLOATING
C2155 VDD.n1266 VSS 0.04fF $ **FLOATING
C2156 VDD.n1267 VSS 0.01fF $ **FLOATING
C2157 VDD.n1268 VSS 0.00fF $ **FLOATING
C2158 VDD.n1269 VSS 0.01fF $ **FLOATING
C2159 VDD.n1270 VSS 0.01fF $ **FLOATING
C2160 VDD.n1271 VSS 0.03fF $ **FLOATING
C2161 VDD.n1272 VSS 0.09fF $ **FLOATING
C2162 VDD.n1273 VSS 0.01fF $ **FLOATING
C2163 VDD.n1274 VSS 4.15fF $ **FLOATING
C2164 VDD.n1276 VSS 0.01fF $ **FLOATING
C2165 VDD.n1277 VSS 0.03fF $ **FLOATING
C2166 VDD.n1278 VSS 0.04fF $ **FLOATING
C2167 VDD.n1279 VSS 0.01fF $ **FLOATING
C2168 VDD.n1280 VSS 0.00fF $ **FLOATING
C2169 VDD.n1281 VSS 0.01fF $ **FLOATING
C2170 VDD.n1282 VSS 0.01fF $ **FLOATING
C2171 VDD.n1283 VSS 0.03fF $ **FLOATING
C2172 VDD.n1284 VSS 0.09fF $ **FLOATING
C2173 VDD.n1285 VSS 0.00fF $ **FLOATING
C2174 VDD.n1286 VSS 0.01fF $ **FLOATING
C2175 VDD.n1287 VSS 0.03fF $ **FLOATING
C2176 VDD.n1288 VSS 0.04fF $ **FLOATING
C2177 VDD.n1289 VSS 0.07fF $ **FLOATING
C2178 VDD.n1290 VSS 0.00fF $ **FLOATING
C2179 VDD.n1291 VSS 0.01fF $ **FLOATING
C2180 VDD.n1292 VSS 0.03fF $ **FLOATING
C2181 VDD.n1293 VSS 0.04fF $ **FLOATING
C2182 VDD.n1294 VSS 0.07fF $ **FLOATING
C2183 VDD.n1295 VSS 0.00fF $ **FLOATING
C2184 VDD.n1296 VSS 0.01fF $ **FLOATING
C2185 VDD.n1297 VSS 0.00fF $ **FLOATING
C2186 VDD.n1298 VSS 0.01fF $ **FLOATING
C2187 VDD.n1299 VSS 0.01fF $ **FLOATING
C2188 VDD.n1300 VSS 0.02fF $ **FLOATING
C2189 VDD.n1301 VSS 0.01fF $ **FLOATING
C2190 VDD.n1302 VSS 8.92fF $ **FLOATING
C2191 VDD.n1303 VSS 0.06fF $ **FLOATING
C2192 VDD.n1304 VSS 0.13fF $ **FLOATING
C2193 VDD.n1305 VSS 5.73fF $ **FLOATING
C2194 VDD.n1306 VSS 0.07fF $ **FLOATING
C2195 VDD.n1307 VSS 0.05fF $ **FLOATING
C2196 VDD.n1308 VSS 0.13fF $ **FLOATING
C2197 VDD.n1309 VSS 0.05fF $ **FLOATING
C2198 VDD.n1310 VSS 0.13fF $ **FLOATING
C2199 VDD.n1311 VSS 0.06fF $ **FLOATING
C2200 VDD.n1312 VSS 0.13fF $ **FLOATING
C2201 VDD.n1313 VSS 0.05fF $ **FLOATING
C2202 VDD.n1314 VSS 0.13fF $ **FLOATING
C2203 VDD.n1315 VSS 5.73fF $ **FLOATING
C2204 VDD.n1316 VSS 0.07fF $ **FLOATING
C2205 VDD.n1317 VSS 0.04fF $ **FLOATING
C2206 VDD.n1318 VSS 0.13fF $ **FLOATING
C2207 VDD.n1319 VSS 0.06fF $ **FLOATING
C2208 VDD.n1320 VSS 0.13fF $ **FLOATING
C2209 VDD.n1321 VSS 0.06fF $ **FLOATING
C2210 VDD.n1322 VSS 0.13fF $ **FLOATING
C2211 VDD.n1323 VSS 5.73fF $ **FLOATING
C2212 VDD.n1324 VSS 0.06fF $ **FLOATING
C2213 VDD.n1325 VSS 0.05fF $ **FLOATING
C2214 VDD.n1326 VSS 0.13fF $ **FLOATING
C2215 VDD.n1327 VSS 0.06fF $ **FLOATING
C2216 VDD.n1328 VSS 0.13fF $ **FLOATING
C2217 VDD.n1329 VSS 0.06fF $ **FLOATING
C2218 VDD.n1330 VSS 0.13fF $ **FLOATING
C2219 VDD.n1331 VSS 5.73fF $ **FLOATING
C2220 VDD.n1332 VSS 0.06fF $ **FLOATING
C2221 VDD.n1333 VSS 0.05fF $ **FLOATING
C2222 VDD.n1334 VSS 0.13fF $ **FLOATING
C2223 VDD.n1335 VSS 0.06fF $ **FLOATING
C2224 VDD.n1336 VSS 0.13fF $ **FLOATING
C2225 VDD.n1337 VSS 0.06fF $ **FLOATING
C2226 VDD.n1338 VSS 0.13fF $ **FLOATING
C2227 VDD.n1339 VSS 5.73fF $ **FLOATING
C2228 VDD.n1340 VSS 0.07fF $ **FLOATING
C2229 VDD.n1341 VSS 0.05fF $ **FLOATING
C2230 VDD.n1342 VSS 0.13fF $ **FLOATING
C2231 VDD.n1343 VSS 0.05fF $ **FLOATING
C2232 VDD.n1344 VSS 0.13fF $ **FLOATING
C2233 VDD.n1345 VSS 0.06fF $ **FLOATING
C2234 VDD.n1346 VSS 0.13fF $ **FLOATING
C2235 VDD.n1347 VSS 0.05fF $ **FLOATING
C2236 VDD.n1348 VSS 0.13fF $ **FLOATING
C2237 VDD.n1349 VSS 5.73fF $ **FLOATING
C2238 VDD.n1350 VSS 0.07fF $ **FLOATING
C2239 VDD.n1351 VSS 0.04fF $ **FLOATING
C2240 VDD.n1352 VSS 0.13fF $ **FLOATING
C2241 VDD.n1353 VSS 0.06fF $ **FLOATING
C2242 VDD.n1354 VSS 0.13fF $ **FLOATING
C2243 VDD.n1355 VSS 0.06fF $ **FLOATING
C2244 VDD.n1356 VSS 0.13fF $ **FLOATING
C2245 VDD.n1357 VSS 5.73fF $ **FLOATING
C2246 VDD.n1358 VSS 0.06fF $ **FLOATING
C2247 VDD.n1359 VSS 0.05fF $ **FLOATING
C2248 VDD.n1360 VSS 0.13fF $ **FLOATING
C2249 VDD.n1361 VSS 0.06fF $ **FLOATING
C2250 VDD.n1362 VSS 0.13fF $ **FLOATING
C2251 VDD.n1363 VSS 0.06fF $ **FLOATING
C2252 VDD.n1364 VSS 0.13fF $ **FLOATING
C2253 VDD.n1365 VSS 5.73fF $ **FLOATING
C2254 VDD.n1366 VSS 0.06fF $ **FLOATING
C2255 VDD.n1367 VSS 0.05fF $ **FLOATING
C2256 VDD.n1368 VSS 0.13fF $ **FLOATING
C2257 VDD.n1369 VSS 0.06fF $ **FLOATING
C2258 VDD.n1370 VSS 0.13fF $ **FLOATING
C2259 VDD.n1371 VSS 0.06fF $ **FLOATING
C2260 VDD.n1372 VSS 0.13fF $ **FLOATING
C2261 VDD.n1373 VSS 5.73fF $ **FLOATING
C2262 VDD.n1374 VSS 0.07fF $ **FLOATING
C2263 VDD.n1375 VSS 0.05fF $ **FLOATING
C2264 VDD.n1376 VSS 0.13fF $ **FLOATING
C2265 VDD.n1377 VSS 0.05fF $ **FLOATING
C2266 VDD.n1378 VSS 0.13fF $ **FLOATING
C2267 VDD.n1379 VSS 0.06fF $ **FLOATING
C2268 VDD.n1380 VSS 0.13fF $ **FLOATING
C2269 VDD.n1381 VSS 0.05fF $ **FLOATING
C2270 VDD.n1382 VSS 0.13fF $ **FLOATING
C2271 VDD.n1383 VSS 5.73fF $ **FLOATING
C2272 VDD.n1384 VSS 0.07fF $ **FLOATING
C2273 VDD.n1385 VSS 0.04fF $ **FLOATING
C2274 VDD.n1386 VSS 0.13fF $ **FLOATING
C2275 VDD.n1387 VSS 0.06fF $ **FLOATING
C2276 VDD.n1388 VSS 0.13fF $ **FLOATING
C2277 VDD.n1389 VSS 0.06fF $ **FLOATING
C2278 VDD.n1390 VSS 0.13fF $ **FLOATING
C2279 VDD.n1391 VSS 5.73fF $ **FLOATING
C2280 VDD.n1392 VSS 0.06fF $ **FLOATING
C2281 VDD.n1393 VSS 0.05fF $ **FLOATING
C2282 VDD.n1394 VSS 0.13fF $ **FLOATING
C2283 VDD.n1395 VSS 0.06fF $ **FLOATING
C2284 VDD.n1396 VSS 0.13fF $ **FLOATING
C2285 VDD.n1397 VSS 0.06fF $ **FLOATING
C2286 VDD.n1398 VSS 0.13fF $ **FLOATING
C2287 VDD.n1399 VSS 5.73fF $ **FLOATING
C2288 VDD.n1400 VSS 0.06fF $ **FLOATING
C2289 VDD.n1401 VSS 0.05fF $ **FLOATING
C2290 VDD.n1402 VSS 0.13fF $ **FLOATING
C2291 VDD.n1403 VSS 0.06fF $ **FLOATING
C2292 VDD.n1404 VSS 0.13fF $ **FLOATING
C2293 VDD.n1405 VSS 0.06fF $ **FLOATING
C2294 VDD.n1406 VSS 0.13fF $ **FLOATING
C2295 VDD.n1407 VSS 5.73fF $ **FLOATING
C2296 VDD.n1408 VSS 0.07fF $ **FLOATING
C2297 VDD.n1409 VSS 0.05fF $ **FLOATING
C2298 VDD.n1410 VSS 0.13fF $ **FLOATING
C2299 VDD.n1411 VSS 0.05fF $ **FLOATING
C2300 VDD.n1412 VSS 0.13fF $ **FLOATING
C2301 VDD.n1413 VSS 0.06fF $ **FLOATING
C2302 VDD.n1414 VSS 0.13fF $ **FLOATING
C2303 VDD.n1415 VSS 0.05fF $ **FLOATING
C2304 VDD.n1416 VSS 0.13fF $ **FLOATING
C2305 VDD.n1417 VSS 7.91fF $ **FLOATING
C2306 VDD.n1418 VSS 0.07fF $ **FLOATING
C2307 VDD.n1419 VSS 0.04fF $ **FLOATING
C2308 VDD.n1420 VSS 0.13fF $ **FLOATING
C2309 VDD.n1421 VSS 0.06fF $ **FLOATING
C2310 VDD.n1422 VSS 0.13fF $ **FLOATING
C2311 VDD.n1423 VSS 0.06fF $ **FLOATING
C2312 VDD.n1424 VSS 0.14fF $ **FLOATING
C2313 VDD.n1425 VSS 0.84fF $ **FLOATING
C2314 VDD.n1426 VSS 0.65fF $ **FLOATING
C2315 VDD.n1427 VSS 0.01fF $ **FLOATING
C2316 VDD.n1428 VSS 0.02fF $ **FLOATING
C2317 VDD.n1429 VSS 0.04fF $ **FLOATING
C2318 VDD.n1430 VSS 0.07fF $ **FLOATING
C2319 VDD.n1431 VSS 0.00fF $ **FLOATING
C2320 VDD.n1432 VSS 0.06fF $ **FLOATING
C2321 VDD.n1434 VSS 3.99fF $ **FLOATING
C2322 VDD.n1435 VSS 3.99fF $ **FLOATING
C2323 VDD.n1437 VSS 0.06fF $ **FLOATING
C2324 VDD.n1438 VSS 0.01fF $ **FLOATING
C2325 VDD.n1439 VSS 0.01fF $ **FLOATING
C2326 VDD.n1440 VSS 0.00fF $ **FLOATING
C2327 VDD.n1441 VSS 0.01fF $ **FLOATING
C2328 VDD.n1442 VSS 0.01fF $ **FLOATING
C2329 VDD.n1443 VSS 0.02fF $ **FLOATING
C2330 VDD.n1444 VSS 0.01fF $ **FLOATING
C2331 VDD.n1445 VSS 0.03fF $ **FLOATING
C2332 VDD.n1446 VSS 0.02fF $ **FLOATING
C2333 VDD.n1447 VSS 0.01fF $ **FLOATING
C2334 VDD.n1448 VSS 1.05fF $ **FLOATING
C2335 VDD.n1449 VSS 0.03fF $ **FLOATING
C2336 VDD.n1450 VSS 3.24fF $ **FLOATING
C2337 VDD.n1451 VSS 0.01fF $ **FLOATING
C2338 VDD.n1452 VSS 0.00fF $ **FLOATING
C2339 VDD.n1453 VSS 0.01fF $ **FLOATING
C2340 VDD.n1454 VSS 0.01fF $ **FLOATING
C2341 VDD.n1455 VSS 0.06fF $ **FLOATING
C2342 VDD.n1456 VSS 0.01fF $ **FLOATING
C2343 VDD.n1457 VSS 0.07fF $ **FLOATING
C2344 VDD.n1458 VSS 0.01fF $ **FLOATING
C2345 VDD.n1459 VSS 0.07fF $ **FLOATING
C2346 VDD.n1460 VSS 0.03fF $ **FLOATING
C2347 VDD.n1461 VSS 0.03fF $ **FLOATING
C2348 VDD.n1462 VSS 0.03fF $ **FLOATING
C2349 VDD.n1463 VSS 0.01fF $ **FLOATING
C2350 VDD.n1464 VSS 0.00fF $ **FLOATING
C2351 VDD.n1465 VSS 0.01fF $ **FLOATING
C2352 VDD.n1466 VSS 0.01fF $ **FLOATING
C2353 VDD.n1467 VSS 0.09fF $ **FLOATING
C2354 VDD.n1468 VSS 0.01fF $ **FLOATING
C2355 VDD.n1469 VSS 0.07fF $ **FLOATING
C2356 VDD.n1470 VSS 0.01fF $ **FLOATING
C2357 VDD.n1471 VSS 0.07fF $ **FLOATING
C2358 VDD.n1472 VSS 0.01fF $ **FLOATING
C2359 VDD.n1473 VSS 0.04fF $ **FLOATING
C2360 VDD.n1474 VSS 0.01fF $ **FLOATING
C2361 VDD.n1475 VSS 0.04fF $ **FLOATING
C2362 VDD.n1476 VSS 0.00fF $ **FLOATING
C2363 VDD.n1477 VSS 0.06fF $ **FLOATING
C2364 VDD.n1479 VSS 3.99fF $ **FLOATING
C2365 VDD.n1480 VSS 3.99fF $ **FLOATING
C2366 VDD.n1482 VSS 0.06fF $ **FLOATING
C2367 VDD.n1483 VSS 0.13fF $ **FLOATING
C2368 VDD.n1484 VSS 5.73fF $ **FLOATING
C2369 VDD.n1485 VSS 0.06fF $ **FLOATING
C2370 VDD.n1486 VSS 0.05fF $ **FLOATING
C2371 VDD.n1487 VSS 0.13fF $ **FLOATING
C2372 VDD.n1488 VSS 0.06fF $ **FLOATING
C2373 VDD.n1489 VSS 0.13fF $ **FLOATING
C2374 VDD.n1490 VSS 0.06fF $ **FLOATING
C2375 VDD.n1491 VSS 0.13fF $ **FLOATING
C2376 VDD.n1492 VSS 5.73fF $ **FLOATING
C2377 VDD.n1493 VSS 0.06fF $ **FLOATING
C2378 VDD.n1494 VSS 0.05fF $ **FLOATING
C2379 VDD.n1495 VSS 0.13fF $ **FLOATING
C2380 VDD.n1496 VSS 0.06fF $ **FLOATING
C2381 VDD.n1497 VSS 0.13fF $ **FLOATING
C2382 VDD.n1498 VSS 0.06fF $ **FLOATING
C2383 VDD.n1499 VSS 0.13fF $ **FLOATING
C2384 VDD.n1500 VSS 5.73fF $ **FLOATING
C2385 VDD.n1501 VSS 0.07fF $ **FLOATING
C2386 VDD.n1502 VSS 0.04fF $ **FLOATING
C2387 VDD.n1503 VSS 0.13fF $ **FLOATING
C2388 VDD.n1504 VSS 0.05fF $ **FLOATING
C2389 VDD.n1505 VSS 0.09fF $ **FLOATING
C2390 VDD.n1506 VSS 9.73fF $ **FLOATING
C2391 VDD.n1507 VSS 0.06fF $ **FLOATING
C2392 VDD.n1508 VSS 0.11fF $ **FLOATING
C2393 VDD.n1509 VSS 0.05fF $ **FLOATING
C2394 VDD.n1510 VSS 0.13fF $ **FLOATING
C2395 VDD.n1511 VSS 5.73fF $ **FLOATING
C2396 VDD.n1512 VSS 0.07fF $ **FLOATING
C2397 VDD.n1513 VSS 0.05fF $ **FLOATING
C2398 VDD.n1514 VSS 0.13fF $ **FLOATING
C2399 VDD.n1515 VSS 0.06fF $ **FLOATING
C2400 VDD.n1516 VSS 0.13fF $ **FLOATING
C2401 VDD.n1517 VSS 0.06fF $ **FLOATING
C2402 VDD.n1518 VSS 0.13fF $ **FLOATING
C2403 VDD.n1519 VSS 7.60fF $ **FLOATING
C2404 VDD.n1520 VSS 0.06fF $ **FLOATING
C2405 VDD.n1521 VSS 0.05fF $ **FLOATING
C2406 VDD.n1522 VSS 0.13fF $ **FLOATING
C2407 VDD.n1523 VSS 0.06fF $ **FLOATING
C2408 VDD.n1524 VSS 0.13fF $ **FLOATING
C2409 VDD.n1525 VSS 0.36fF $ **FLOATING
C2410 VDD.n1526 VSS 0.10fF $ **FLOATING
C2411 VDD.n1527 VSS 2.81fF $ **FLOATING
C2412 VDD.n1528 VSS 0.03fF $ **FLOATING
C2413 VDD.n1529 VSS 2.74fF $ **FLOATING
C2414 VDD.n1530 VSS 0.01fF $ **FLOATING
C2415 VDD.n1531 VSS 0.00fF $ **FLOATING
C2416 VDD.n1532 VSS 0.01fF $ **FLOATING
C2417 VDD.n1533 VSS 0.01fF $ **FLOATING
C2418 VDD.n1534 VSS 0.06fF $ **FLOATING
C2419 VDD.n1535 VSS 0.03fF $ **FLOATING
C2420 VDD.n1536 VSS 0.04fF $ **FLOATING
C2421 VDD.n1537 VSS 0.01fF $ **FLOATING
C2422 VDD.n1538 VSS 0.07fF $ **FLOATING
C2423 VDD.n1539 VSS 0.01fF $ **FLOATING
C2424 VDD.n1540 VSS 0.03fF $ **FLOATING
C2425 VDD.n1541 VSS 0.04fF $ **FLOATING
C2426 VDD.n1542 VSS 0.01fF $ **FLOATING
C2427 VDD.n1543 VSS 0.07fF $ **FLOATING
C2428 VDD.n1544 VSS 0.01fF $ **FLOATING
C2429 VDD.n1545 VSS 0.03fF $ **FLOATING
C2430 VDD.n1546 VSS 0.04fF $ **FLOATING
C2431 VDD.n1547 VSS 0.01fF $ **FLOATING
C2432 VDD.n1548 VSS 0.07fF $ **FLOATING
C2433 VDD.n1549 VSS 0.01fF $ **FLOATING
C2434 VDD.n1550 VSS 0.01fF $ **FLOATING
C2435 VDD.n1551 VSS 0.00fF $ **FLOATING
C2436 VDD.n1552 VSS 0.01fF $ **FLOATING
C2437 VDD.n1553 VSS 0.01fF $ **FLOATING
C2438 VDD.n1554 VSS 0.03fF $ **FLOATING
C2439 VDD.n1555 VSS 0.05fF $ **FLOATING
C2440 VDD.n1556 VSS 0.04fF $ **FLOATING
C2441 VDD.n1557 VSS 0.01fF $ **FLOATING
C2442 VDD.n1558 VSS 0.06fF $ **FLOATING
C2443 VDD.n1560 VSS 4.15fF $ **FLOATING
C2444 VDD.n1561 VSS 62.36fF $ **FLOATING
C2445 vbg.n0 VSS 1.23fF $ **FLOATING
C2446 vbg.n1 VSS 0.03fF $ **FLOATING
C2447 vbg.n2 VSS 0.01fF $ **FLOATING
C2448 vbg.n3 VSS 0.01fF $ **FLOATING
C2449 vbg.n4 VSS 0.00fF $ **FLOATING
C2450 vbg.n5 VSS 0.00fF $ **FLOATING
C2451 vbg.n6 VSS 0.01fF $ **FLOATING
C2452 vbg.n7 VSS 0.01fF $ **FLOATING
C2453 vbg.n8 VSS 0.01fF $ **FLOATING
C2454 vbg.n9 VSS 0.00fF $ **FLOATING
C2455 vbg.n10 VSS 0.01fF $ **FLOATING
C2456 vbg.n11 VSS 0.00fF $ **FLOATING
C2457 vbg.n12 VSS 0.01fF $ **FLOATING
C2458 vbg.n13 VSS 0.00fF $ **FLOATING
C2459 vbg.n14 VSS 0.01fF $ **FLOATING
C2460 vbg.n15 VSS 0.00fF $ **FLOATING
C2461 vbg.n16 VSS 0.00fF $ **FLOATING
C2462 vbg.n17 VSS 0.01fF $ **FLOATING
C2463 vbg.n18 VSS 0.01fF $ **FLOATING
C2464 vbg.n19 VSS 0.01fF $ **FLOATING
C2465 vbg.n20 VSS 0.00fF $ **FLOATING
C2466 vbg.n21 VSS 0.01fF $ **FLOATING
C2467 vbg.n22 VSS 0.00fF $ **FLOATING
C2468 vbg.n23 VSS 0.01fF $ **FLOATING
C2469 vbg.n24 VSS 0.00fF $ **FLOATING
C2470 vbg.n25 VSS 0.01fF $ **FLOATING
C2471 vbg.n26 VSS 0.00fF $ **FLOATING
C2472 vbg.n27 VSS 0.00fF $ **FLOATING
C2473 vbg.n28 VSS 0.01fF $ **FLOATING
C2474 vbg.n29 VSS 0.01fF $ **FLOATING
C2475 vbg.n30 VSS 0.00fF $ **FLOATING
C2476 vbg.n31 VSS 0.00fF $ **FLOATING
C2477 vbg.n32 VSS 0.01fF $ **FLOATING
C2478 vbg.n33 VSS 0.00fF $ **FLOATING
C2479 vbg.n34 VSS 0.01fF $ **FLOATING
C2480 vbg.n35 VSS 0.00fF $ **FLOATING
C2481 vbg.n36 VSS 0.01fF $ **FLOATING
C2482 vbg.n37 VSS 0.00fF $ **FLOATING
C2483 vbg.n38 VSS 0.00fF $ **FLOATING
C2484 vbg.n39 VSS 0.00fF $ **FLOATING
C2485 vbg.n40 VSS 0.01fF $ **FLOATING
C2486 vbg.n41 VSS 0.00fF $ **FLOATING
C2487 vbg.n42 VSS 0.00fF $ **FLOATING
C2488 vbg.n43 VSS 0.01fF $ **FLOATING
C2489 vbg.n44 VSS 0.00fF $ **FLOATING
C2490 vbg.n45 VSS 0.01fF $ **FLOATING
C2491 vbg.n46 VSS 0.00fF $ **FLOATING
C2492 vbg.n47 VSS 0.01fF $ **FLOATING
C2493 vbg.n48 VSS 0.00fF $ **FLOATING
C2494 vbg.n49 VSS 0.00fF $ **FLOATING
C2495 vbg.n50 VSS 0.00fF $ **FLOATING
C2496 vbg.n51 VSS 0.01fF $ **FLOATING
C2497 vbg.n52 VSS 0.00fF $ **FLOATING
C2498 vbg.n53 VSS 0.00fF $ **FLOATING
C2499 vbg.n54 VSS 0.01fF $ **FLOATING
C2500 vbg.n55 VSS 0.00fF $ **FLOATING
C2501 vbg.n56 VSS 0.01fF $ **FLOATING
C2502 vbg.n57 VSS 0.00fF $ **FLOATING
C2503 vbg.n58 VSS 0.01fF $ **FLOATING
C2504 vbg.n59 VSS 0.00fF $ **FLOATING
C2505 vbg.n60 VSS 0.00fF $ **FLOATING
C2506 vbg.n61 VSS 0.00fF $ **FLOATING
C2507 vbg.n62 VSS 0.01fF $ **FLOATING
C2508 vbg.n63 VSS 0.00fF $ **FLOATING
C2509 vbg.n64 VSS 0.00fF $ **FLOATING
C2510 vbg.n65 VSS 0.01fF $ **FLOATING
C2511 vbg.n66 VSS 0.00fF $ **FLOATING
C2512 vbg.n67 VSS 0.01fF $ **FLOATING
C2513 vbg.n68 VSS 0.00fF $ **FLOATING
C2514 vbg.n69 VSS 0.01fF $ **FLOATING
C2515 vbg.n70 VSS 0.00fF $ **FLOATING
C2516 vbg.n71 VSS 0.00fF $ **FLOATING
C2517 vbg.n72 VSS 0.00fF $ **FLOATING
C2518 vbg.n73 VSS 0.01fF $ **FLOATING
C2519 vbg.n74 VSS 0.00fF $ **FLOATING
C2520 vbg.n75 VSS 0.00fF $ **FLOATING
C2521 vbg.n76 VSS 0.01fF $ **FLOATING
C2522 vbg.n77 VSS 0.00fF $ **FLOATING
C2523 vbg.n78 VSS 0.01fF $ **FLOATING
C2524 vbg.n79 VSS 0.00fF $ **FLOATING
C2525 vbg.n80 VSS 0.01fF $ **FLOATING
C2526 vbg.n81 VSS 0.00fF $ **FLOATING
C2527 vbg.n82 VSS 0.00fF $ **FLOATING
C2528 vbg.n83 VSS 0.00fF $ **FLOATING
C2529 vbg.n84 VSS 0.01fF $ **FLOATING
C2530 vbg.n85 VSS 0.01fF $ **FLOATING
C2531 vbg.n86 VSS 0.00fF $ **FLOATING
C2532 vbg.n87 VSS 0.01fF $ **FLOATING
C2533 vbg.n88 VSS 0.00fF $ **FLOATING
C2534 vbg.n89 VSS 0.00fF $ **FLOATING
C2535 vbg.n90 VSS 0.00fF $ **FLOATING
C2536 vbg.n91 VSS 0.00fF $ **FLOATING
C2537 vbg.n92 VSS 0.02fF $ **FLOATING
C2538 vbg.n93 VSS 0.01fF $ **FLOATING
C2539 vbg.n94 VSS 0.00fF $ **FLOATING
C2540 vbg.n95 VSS 0.01fF $ **FLOATING
C2541 vbg.n96 VSS 0.00fF $ **FLOATING
C2542 vbg.n97 VSS 0.01fF $ **FLOATING
C2543 vbg.n98 VSS 0.00fF $ **FLOATING
C2544 vbg.n99 VSS 0.01fF $ **FLOATING
C2545 vbg.n100 VSS 0.00fF $ **FLOATING
C2546 vbg.n101 VSS 0.00fF $ **FLOATING
C2547 vbg.n102 VSS 0.00fF $ **FLOATING
C2548 vbg.n103 VSS 0.00fF $ **FLOATING
C2549 vbg.n104 VSS 0.01fF $ **FLOATING
C2550 vbg.n105 VSS 0.00fF $ **FLOATING
C2551 vbg.n106 VSS 0.01fF $ **FLOATING
C2552 vbg.n107 VSS 0.00fF $ **FLOATING
C2553 vbg.n108 VSS 0.01fF $ **FLOATING
C2554 vbg.n109 VSS 0.00fF $ **FLOATING
C2555 vbg.n110 VSS 0.01fF $ **FLOATING
C2556 vbg.n111 VSS 0.00fF $ **FLOATING
C2557 vbg.n112 VSS 0.00fF $ **FLOATING
C2558 vbg.n113 VSS 0.00fF $ **FLOATING
C2559 vbg.n114 VSS 0.00fF $ **FLOATING
C2560 vbg.n115 VSS 0.01fF $ **FLOATING
C2561 vbg.n116 VSS 0.00fF $ **FLOATING
C2562 vbg.n117 VSS 0.01fF $ **FLOATING
C2563 vbg.n118 VSS 0.00fF $ **FLOATING
C2564 vbg.n119 VSS 0.01fF $ **FLOATING
C2565 vbg.n120 VSS 0.00fF $ **FLOATING
C2566 vbg.n121 VSS 0.01fF $ **FLOATING
C2567 vbg.n122 VSS 0.00fF $ **FLOATING
C2568 vbg.n123 VSS 0.00fF $ **FLOATING
C2569 vbg.n124 VSS 0.00fF $ **FLOATING
C2570 vbg.n125 VSS 0.00fF $ **FLOATING
C2571 vbg.n126 VSS 0.01fF $ **FLOATING
C2572 vbg.n127 VSS 0.00fF $ **FLOATING
C2573 vbg.n128 VSS 0.01fF $ **FLOATING
C2574 vbg.n129 VSS 0.00fF $ **FLOATING
C2575 vbg.n130 VSS 0.01fF $ **FLOATING
C2576 vbg.n131 VSS 0.00fF $ **FLOATING
C2577 vbg.n132 VSS 0.01fF $ **FLOATING
C2578 vbg.n133 VSS 0.00fF $ **FLOATING
C2579 vbg.n134 VSS 0.00fF $ **FLOATING
C2580 vbg.n135 VSS 0.00fF $ **FLOATING
C2581 vbg.n136 VSS 0.00fF $ **FLOATING
C2582 vbg.n137 VSS 0.01fF $ **FLOATING
C2583 vbg.n138 VSS 0.00fF $ **FLOATING
C2584 vbg.n139 VSS 0.01fF $ **FLOATING
C2585 vbg.n140 VSS 0.00fF $ **FLOATING
C2586 vbg.n141 VSS 0.01fF $ **FLOATING
C2587 vbg.n142 VSS 0.01fF $ **FLOATING
C2588 vbg.n143 VSS 0.01fF $ **FLOATING
C2589 vbg.n144 VSS 0.00fF $ **FLOATING
C2590 vbg.n145 VSS 0.00fF $ **FLOATING
C2591 vbg.n146 VSS 0.01fF $ **FLOATING
C2592 vbg.n147 VSS 0.00fF $ **FLOATING
C2593 vbg.n148 VSS 0.01fF $ **FLOATING
C2594 vbg.n149 VSS 0.00fF $ **FLOATING
C2595 vbg.n150 VSS 0.01fF $ **FLOATING
C2596 vbg.n151 VSS 0.00fF $ **FLOATING
C2597 vbg.n152 VSS 0.01fF $ **FLOATING
C2598 vbg.n153 VSS 0.01fF $ **FLOATING
C2599 vbg.n154 VSS 0.01fF $ **FLOATING
C2600 vbg.n155 VSS 0.00fF $ **FLOATING
C2601 vbg.n156 VSS 0.00fF $ **FLOATING
C2602 vbg.n157 VSS 0.01fF $ **FLOATING
C2603 vbg.n158 VSS 0.00fF $ **FLOATING
C2604 vbg.n159 VSS 0.01fF $ **FLOATING
C2605 vbg.n160 VSS 0.00fF $ **FLOATING
C2606 vbg.n161 VSS 0.01fF $ **FLOATING
C2607 vbg.n162 VSS 0.00fF $ **FLOATING
C2608 vbg.n163 VSS 0.01fF $ **FLOATING
C2609 vbg.n164 VSS 0.01fF $ **FLOATING
C2610 vbg.n165 VSS 0.01fF $ **FLOATING
C2611 vbg.n166 VSS 0.00fF $ **FLOATING
C2612 vbg.n167 VSS 0.00fF $ **FLOATING
C2613 vbg.n168 VSS 0.02fF $ **FLOATING
C2614 vbg.n169 VSS 0.01fF $ **FLOATING
C2615 vbg.n170 VSS 0.03fF $ **FLOATING
C2616 vbg.n171 VSS 38.53fF $ **FLOATING
C2617 vbg.n172 VSS 6.97fF $ **FLOATING
C2618 sky130_asc_res_xhigh_po_2p85_1_5/Rin VSS 6.60fF
C2619 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# VSS 2.70fF
C2620 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# VSS 2.70fF
C2621 sky130_asc_res_xhigh_po_2p85_1_3/Rin VSS 3.23fF
C2622 sky130_asc_res_xhigh_po_2p85_1_4/Rin VSS 4.07fF
C2623 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# VSS 2.70fF
C2624 va VSS 162.71fF
C2625 sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# VSS 2.70fF
C2626 sky130_asc_res_xhigh_po_2p85_1_1/Rin VSS 4.40fF
C2627 sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# VSS 2.70fF
C2628 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS 10.35fF
C2629 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS 3.54fF
C2630 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# VSS 2.90fF
C2631 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# VSS 2.70fF
C2632 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS 58.51fF
C2633 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# VSS 2.86fF
C2634 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# VSS 2.70fF
C2635 sky130_asc_res_xhigh_po_2p85_1_17/Rin VSS 3.90fF
C2636 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# VSS 2.70fF
C2637 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# VSS 2.70fF
C2638 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# VSS 2.70fF
C2639 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# VSS 2.70fF
C2640 sky130_asc_res_xhigh_po_2p85_1_15/Rin VSS 5.80fF
C2641 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# VSS 2.86fF
C2642 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# VSS 2.70fF
C2643 sky130_asc_res_xhigh_po_2p85_1_25/Rin VSS 4.29fF
C2644 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# VSS 2.70fF
C2645 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS 14.93fF
C2646 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# VSS 2.70fF
C2647 sky130_asc_res_xhigh_po_2p85_1_24/Rin VSS 5.51fF
C2648 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# VSS 2.70fF
C2649 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# VSS 2.70fF
C2650 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# VSS 2.85fF
C2651 sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# VSS 2.70fF
C2652 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# VSS 2.70fF
C2653 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# VSS 2.70fF
C2654 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# VSS 2.70fF
C2655 sky130_asc_res_xhigh_po_2p85_1_11/Rin VSS 5.36fF
C2656 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# VSS 2.70fF
C2657 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# VSS 2.70fF
C2658 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS 3.06fF
C2659 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# VSS 2.70fF
C2660 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# VSS 2.70fF
C2661 sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# VSS 2.86fF
C2662 sky130_asc_res_xhigh_po_2p85_1_29/Rin VSS 4.48fF
C2663 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# VSS 2.70fF
C2664 sky130_asc_cap_mim_m3_1_4/Cout VSS 130.29fF
C2665 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# VSS 2.70fF
C2666 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# VSS 2.70fF
C2667 sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# VSS 2.70fF

**** begin user architecture code

.lib /farmshare/home/classes/ee/272/PDKs/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.option savecurrents
.param R3val='22.187k'
.param alpha='1'
.param R2R3ratio='5.6555038*alpha'
.param R2val='R3val*R2R3ratio'
.param R4R2ratio='0.79694273'
.param R4val='R2val*R4R2ratio'
.nodeset v(vgate)=1.4
.param VDD=1.8
.control
save all  @m.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm5.msky130_fd_pr__nfet_01v8_lvt[gm]  @m.xm6.msky130_fd_pr__nfet_01v8_lvt[gm]  @m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]  @m.xm8.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm9.msky130_fd_pr__nfet_01v8_lvt[gm]  @m.xm13.msky130_fd_pr__pfet_01v8_lvt[gm]

op

let id8=@m.xm8.msky130_fd_pr__pfet_01v8_lvt[id]
let id1=@m.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
let vth5=@m.xm5.msky130_fd_pr__nfet_01v8_lvt[vth]
let vth6=@m.xm6.msky130_fd_pr__nfet_01v8_lvt[vth]
let wm8=@m.xm8.msky130_fd_pr__pfet_01v8_lvt[w]
let mm8=@m.xm8.msky130_fd_pr__pfet_01v8_lvt[m]
let weff8=wm8*mm8
let jd8=id8/weff8
let wm1=@m.xm1.msky130_fd_pr__pfet_01v8_lvt[w]
let mm1=@m.xm1.msky130_fd_pr__pfet_01v8_lvt[m]
let weff1=wm1*mm1
let jd1=id1/weff1
let wm13=@m.xm13.msky130_fd_pr__pfet_01v8_lvt[w]
let mm13=@m.xm13.msky130_fd_pr__pfet_01v8_lvt[m]
let weff13=wm13*mm13
let id13=@m.xm13.msky130_fd_pr__pfet_01v8_lvt[id]
let jd13=id13/weff13
let gm13=@m.xm13.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm3=@m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm4=@m.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm5=@m.xm5.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm6=@m.xm6.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm7=@m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm8=@m.xm8.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm9=@m.xm9.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm1=@m.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm2=@m.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
let vdsat1=2/(gm1/vm1#branch)
let vdsat2=2/(gm2/vm2#branch)
let vdsat3=2/(gm3/vm3#branch)
let vdsat4=2/(gm4/@m.xm4.msky130_fd_pr__pfet_01v8_lvt[id])
let vdsat5=2/(gm5/@m.xm5.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat6=2/(gm6/@m.xm6.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat7=2/(gm7/@m.xm7.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat8=2/(gm8/@m.xm8.msky130_fd_pr__pfet_01v8_lvt[id])
let vdsat9=2/(gm9/@m.xm9.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat13=2/(gm13/@m.xm13.msky130_fd_pr__pfet_01v8_lvt[id])

write 
print vbg vgate vg va vb vx vq
print vdsat1 vdsat2 vdsat3 vdsat4   vdsat5 vdsat6 vdsat7 vdsat8 vdsat9 vdsat13 
unset askquit
quit
.endc


**** end user architecture code
**.ends
.GLOBAL VDD 
.GLOBAL GND 
** flattened .save nodes
.save I(Vr4)
.save I(Vr2)
.save I(Vm1)
.save I(Vm2)
.save I(Vm3)
.save I(Vr1)
.save I(Vq2)
.end 
