VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.330 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 3.880 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 3.880 8.650 ;
        RECT 3.465 8.245 3.635 8.450 ;
        RECT 3.465 8.130 3.640 8.245 ;
        RECT 3.470 1.755 3.640 8.130 ;
      LAYER mcon ;
        RECT 3.470 1.835 3.640 8.165 ;
      LAYER met1 ;
        RECT 3.440 1.775 3.670 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 1.180 1.870 1.350 8.245 ;
        RECT 1.175 1.755 1.350 1.870 ;
        RECT 1.175 1.350 1.345 1.755 ;
        RECT 0.940 1.050 3.880 1.350 ;
      LAYER mcon ;
        RECT 1.180 1.835 1.350 8.165 ;
      LAYER met1 ;
        RECT 1.150 1.775 1.380 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 1.470 3.880 9.700 ;
        RECT 0.940 1.465 3.880 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 3.880 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 3.880 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 3.880 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 3.880 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1
END LIBRARY

