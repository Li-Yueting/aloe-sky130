VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 53.600 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.965 5.085 6.435 ;
        RECT 8.315 2.965 11.785 6.435 ;
        RECT 15.015 2.965 18.485 6.435 ;
        RECT 21.715 2.965 25.185 6.435 ;
        RECT 28.415 2.965 31.885 6.435 ;
        RECT 35.115 2.965 38.585 6.435 ;
        RECT 41.815 2.965 45.285 6.435 ;
        RECT 48.515 2.965 51.985 6.435 ;
      LAYER mcon ;
        RECT 1.980 5.830 2.150 6.000 ;
        RECT 2.480 5.830 2.650 6.000 ;
        RECT 2.980 5.830 3.150 6.000 ;
        RECT 3.480 5.830 3.650 6.000 ;
        RECT 3.980 5.830 4.150 6.000 ;
        RECT 4.480 5.830 4.650 6.000 ;
        RECT 1.980 5.330 2.150 5.500 ;
        RECT 2.480 5.330 2.650 5.500 ;
        RECT 2.980 5.330 3.150 5.500 ;
        RECT 3.480 5.330 3.650 5.500 ;
        RECT 3.980 5.330 4.150 5.500 ;
        RECT 4.480 5.330 4.650 5.500 ;
        RECT 1.980 4.830 2.150 5.000 ;
        RECT 2.480 4.830 2.650 5.000 ;
        RECT 2.980 4.830 3.150 5.000 ;
        RECT 3.480 4.830 3.650 5.000 ;
        RECT 3.980 4.830 4.150 5.000 ;
        RECT 4.480 4.830 4.650 5.000 ;
        RECT 1.980 4.330 2.150 4.500 ;
        RECT 2.480 4.330 2.650 4.500 ;
        RECT 2.980 4.330 3.150 4.500 ;
        RECT 3.480 4.330 3.650 4.500 ;
        RECT 3.980 4.330 4.150 4.500 ;
        RECT 4.480 4.330 4.650 4.500 ;
        RECT 1.980 3.830 2.150 4.000 ;
        RECT 2.480 3.830 2.650 4.000 ;
        RECT 2.980 3.830 3.150 4.000 ;
        RECT 3.480 3.830 3.650 4.000 ;
        RECT 3.980 3.830 4.150 4.000 ;
        RECT 4.480 3.830 4.650 4.000 ;
        RECT 1.980 3.330 2.150 3.500 ;
        RECT 2.480 3.330 2.650 3.500 ;
        RECT 2.980 3.330 3.150 3.500 ;
        RECT 3.480 3.330 3.650 3.500 ;
        RECT 3.980 3.330 4.150 3.500 ;
        RECT 4.480 3.330 4.650 3.500 ;
        RECT 8.680 5.830 8.850 6.000 ;
        RECT 9.180 5.830 9.350 6.000 ;
        RECT 9.680 5.830 9.850 6.000 ;
        RECT 10.180 5.830 10.350 6.000 ;
        RECT 10.680 5.830 10.850 6.000 ;
        RECT 11.180 5.830 11.350 6.000 ;
        RECT 8.680 5.330 8.850 5.500 ;
        RECT 9.180 5.330 9.350 5.500 ;
        RECT 9.680 5.330 9.850 5.500 ;
        RECT 10.180 5.330 10.350 5.500 ;
        RECT 10.680 5.330 10.850 5.500 ;
        RECT 11.180 5.330 11.350 5.500 ;
        RECT 8.680 4.830 8.850 5.000 ;
        RECT 9.180 4.830 9.350 5.000 ;
        RECT 9.680 4.830 9.850 5.000 ;
        RECT 10.180 4.830 10.350 5.000 ;
        RECT 10.680 4.830 10.850 5.000 ;
        RECT 11.180 4.830 11.350 5.000 ;
        RECT 8.680 4.330 8.850 4.500 ;
        RECT 9.180 4.330 9.350 4.500 ;
        RECT 9.680 4.330 9.850 4.500 ;
        RECT 10.180 4.330 10.350 4.500 ;
        RECT 10.680 4.330 10.850 4.500 ;
        RECT 11.180 4.330 11.350 4.500 ;
        RECT 8.680 3.830 8.850 4.000 ;
        RECT 9.180 3.830 9.350 4.000 ;
        RECT 9.680 3.830 9.850 4.000 ;
        RECT 10.180 3.830 10.350 4.000 ;
        RECT 10.680 3.830 10.850 4.000 ;
        RECT 11.180 3.830 11.350 4.000 ;
        RECT 8.680 3.330 8.850 3.500 ;
        RECT 9.180 3.330 9.350 3.500 ;
        RECT 9.680 3.330 9.850 3.500 ;
        RECT 10.180 3.330 10.350 3.500 ;
        RECT 10.680 3.330 10.850 3.500 ;
        RECT 11.180 3.330 11.350 3.500 ;
        RECT 15.380 5.830 15.550 6.000 ;
        RECT 15.880 5.830 16.050 6.000 ;
        RECT 16.380 5.830 16.550 6.000 ;
        RECT 16.880 5.830 17.050 6.000 ;
        RECT 17.380 5.830 17.550 6.000 ;
        RECT 17.880 5.830 18.050 6.000 ;
        RECT 15.380 5.330 15.550 5.500 ;
        RECT 15.880 5.330 16.050 5.500 ;
        RECT 16.380 5.330 16.550 5.500 ;
        RECT 16.880 5.330 17.050 5.500 ;
        RECT 17.380 5.330 17.550 5.500 ;
        RECT 17.880 5.330 18.050 5.500 ;
        RECT 15.380 4.830 15.550 5.000 ;
        RECT 15.880 4.830 16.050 5.000 ;
        RECT 16.380 4.830 16.550 5.000 ;
        RECT 16.880 4.830 17.050 5.000 ;
        RECT 17.380 4.830 17.550 5.000 ;
        RECT 17.880 4.830 18.050 5.000 ;
        RECT 15.380 4.330 15.550 4.500 ;
        RECT 15.880 4.330 16.050 4.500 ;
        RECT 16.380 4.330 16.550 4.500 ;
        RECT 16.880 4.330 17.050 4.500 ;
        RECT 17.380 4.330 17.550 4.500 ;
        RECT 17.880 4.330 18.050 4.500 ;
        RECT 15.380 3.830 15.550 4.000 ;
        RECT 15.880 3.830 16.050 4.000 ;
        RECT 16.380 3.830 16.550 4.000 ;
        RECT 16.880 3.830 17.050 4.000 ;
        RECT 17.380 3.830 17.550 4.000 ;
        RECT 17.880 3.830 18.050 4.000 ;
        RECT 15.380 3.330 15.550 3.500 ;
        RECT 15.880 3.330 16.050 3.500 ;
        RECT 16.380 3.330 16.550 3.500 ;
        RECT 16.880 3.330 17.050 3.500 ;
        RECT 17.380 3.330 17.550 3.500 ;
        RECT 17.880 3.330 18.050 3.500 ;
        RECT 22.080 5.830 22.250 6.000 ;
        RECT 22.580 5.830 22.750 6.000 ;
        RECT 23.080 5.830 23.250 6.000 ;
        RECT 23.580 5.830 23.750 6.000 ;
        RECT 24.080 5.830 24.250 6.000 ;
        RECT 24.580 5.830 24.750 6.000 ;
        RECT 22.080 5.330 22.250 5.500 ;
        RECT 22.580 5.330 22.750 5.500 ;
        RECT 23.080 5.330 23.250 5.500 ;
        RECT 23.580 5.330 23.750 5.500 ;
        RECT 24.080 5.330 24.250 5.500 ;
        RECT 24.580 5.330 24.750 5.500 ;
        RECT 22.080 4.830 22.250 5.000 ;
        RECT 22.580 4.830 22.750 5.000 ;
        RECT 23.080 4.830 23.250 5.000 ;
        RECT 23.580 4.830 23.750 5.000 ;
        RECT 24.080 4.830 24.250 5.000 ;
        RECT 24.580 4.830 24.750 5.000 ;
        RECT 22.080 4.330 22.250 4.500 ;
        RECT 22.580 4.330 22.750 4.500 ;
        RECT 23.080 4.330 23.250 4.500 ;
        RECT 23.580 4.330 23.750 4.500 ;
        RECT 24.080 4.330 24.250 4.500 ;
        RECT 24.580 4.330 24.750 4.500 ;
        RECT 22.080 3.830 22.250 4.000 ;
        RECT 22.580 3.830 22.750 4.000 ;
        RECT 23.080 3.830 23.250 4.000 ;
        RECT 23.580 3.830 23.750 4.000 ;
        RECT 24.080 3.830 24.250 4.000 ;
        RECT 24.580 3.830 24.750 4.000 ;
        RECT 22.080 3.330 22.250 3.500 ;
        RECT 22.580 3.330 22.750 3.500 ;
        RECT 23.080 3.330 23.250 3.500 ;
        RECT 23.580 3.330 23.750 3.500 ;
        RECT 24.080 3.330 24.250 3.500 ;
        RECT 24.580 3.330 24.750 3.500 ;
        RECT 28.780 5.830 28.950 6.000 ;
        RECT 29.280 5.830 29.450 6.000 ;
        RECT 29.780 5.830 29.950 6.000 ;
        RECT 30.280 5.830 30.450 6.000 ;
        RECT 30.780 5.830 30.950 6.000 ;
        RECT 31.280 5.830 31.450 6.000 ;
        RECT 28.780 5.330 28.950 5.500 ;
        RECT 29.280 5.330 29.450 5.500 ;
        RECT 29.780 5.330 29.950 5.500 ;
        RECT 30.280 5.330 30.450 5.500 ;
        RECT 30.780 5.330 30.950 5.500 ;
        RECT 31.280 5.330 31.450 5.500 ;
        RECT 28.780 4.830 28.950 5.000 ;
        RECT 29.280 4.830 29.450 5.000 ;
        RECT 29.780 4.830 29.950 5.000 ;
        RECT 30.280 4.830 30.450 5.000 ;
        RECT 30.780 4.830 30.950 5.000 ;
        RECT 31.280 4.830 31.450 5.000 ;
        RECT 28.780 4.330 28.950 4.500 ;
        RECT 29.280 4.330 29.450 4.500 ;
        RECT 29.780 4.330 29.950 4.500 ;
        RECT 30.280 4.330 30.450 4.500 ;
        RECT 30.780 4.330 30.950 4.500 ;
        RECT 31.280 4.330 31.450 4.500 ;
        RECT 28.780 3.830 28.950 4.000 ;
        RECT 29.280 3.830 29.450 4.000 ;
        RECT 29.780 3.830 29.950 4.000 ;
        RECT 30.280 3.830 30.450 4.000 ;
        RECT 30.780 3.830 30.950 4.000 ;
        RECT 31.280 3.830 31.450 4.000 ;
        RECT 28.780 3.330 28.950 3.500 ;
        RECT 29.280 3.330 29.450 3.500 ;
        RECT 29.780 3.330 29.950 3.500 ;
        RECT 30.280 3.330 30.450 3.500 ;
        RECT 30.780 3.330 30.950 3.500 ;
        RECT 31.280 3.330 31.450 3.500 ;
        RECT 35.480 5.830 35.650 6.000 ;
        RECT 35.980 5.830 36.150 6.000 ;
        RECT 36.480 5.830 36.650 6.000 ;
        RECT 36.980 5.830 37.150 6.000 ;
        RECT 37.480 5.830 37.650 6.000 ;
        RECT 37.980 5.830 38.150 6.000 ;
        RECT 35.480 5.330 35.650 5.500 ;
        RECT 35.980 5.330 36.150 5.500 ;
        RECT 36.480 5.330 36.650 5.500 ;
        RECT 36.980 5.330 37.150 5.500 ;
        RECT 37.480 5.330 37.650 5.500 ;
        RECT 37.980 5.330 38.150 5.500 ;
        RECT 35.480 4.830 35.650 5.000 ;
        RECT 35.980 4.830 36.150 5.000 ;
        RECT 36.480 4.830 36.650 5.000 ;
        RECT 36.980 4.830 37.150 5.000 ;
        RECT 37.480 4.830 37.650 5.000 ;
        RECT 37.980 4.830 38.150 5.000 ;
        RECT 35.480 4.330 35.650 4.500 ;
        RECT 35.980 4.330 36.150 4.500 ;
        RECT 36.480 4.330 36.650 4.500 ;
        RECT 36.980 4.330 37.150 4.500 ;
        RECT 37.480 4.330 37.650 4.500 ;
        RECT 37.980 4.330 38.150 4.500 ;
        RECT 35.480 3.830 35.650 4.000 ;
        RECT 35.980 3.830 36.150 4.000 ;
        RECT 36.480 3.830 36.650 4.000 ;
        RECT 36.980 3.830 37.150 4.000 ;
        RECT 37.480 3.830 37.650 4.000 ;
        RECT 37.980 3.830 38.150 4.000 ;
        RECT 35.480 3.330 35.650 3.500 ;
        RECT 35.980 3.330 36.150 3.500 ;
        RECT 36.480 3.330 36.650 3.500 ;
        RECT 36.980 3.330 37.150 3.500 ;
        RECT 37.480 3.330 37.650 3.500 ;
        RECT 37.980 3.330 38.150 3.500 ;
        RECT 42.180 5.830 42.350 6.000 ;
        RECT 42.680 5.830 42.850 6.000 ;
        RECT 43.180 5.830 43.350 6.000 ;
        RECT 43.680 5.830 43.850 6.000 ;
        RECT 44.180 5.830 44.350 6.000 ;
        RECT 44.680 5.830 44.850 6.000 ;
        RECT 42.180 5.330 42.350 5.500 ;
        RECT 42.680 5.330 42.850 5.500 ;
        RECT 43.180 5.330 43.350 5.500 ;
        RECT 43.680 5.330 43.850 5.500 ;
        RECT 44.180 5.330 44.350 5.500 ;
        RECT 44.680 5.330 44.850 5.500 ;
        RECT 42.180 4.830 42.350 5.000 ;
        RECT 42.680 4.830 42.850 5.000 ;
        RECT 43.180 4.830 43.350 5.000 ;
        RECT 43.680 4.830 43.850 5.000 ;
        RECT 44.180 4.830 44.350 5.000 ;
        RECT 44.680 4.830 44.850 5.000 ;
        RECT 42.180 4.330 42.350 4.500 ;
        RECT 42.680 4.330 42.850 4.500 ;
        RECT 43.180 4.330 43.350 4.500 ;
        RECT 43.680 4.330 43.850 4.500 ;
        RECT 44.180 4.330 44.350 4.500 ;
        RECT 44.680 4.330 44.850 4.500 ;
        RECT 42.180 3.830 42.350 4.000 ;
        RECT 42.680 3.830 42.850 4.000 ;
        RECT 43.180 3.830 43.350 4.000 ;
        RECT 43.680 3.830 43.850 4.000 ;
        RECT 44.180 3.830 44.350 4.000 ;
        RECT 44.680 3.830 44.850 4.000 ;
        RECT 42.180 3.330 42.350 3.500 ;
        RECT 42.680 3.330 42.850 3.500 ;
        RECT 43.180 3.330 43.350 3.500 ;
        RECT 43.680 3.330 43.850 3.500 ;
        RECT 44.180 3.330 44.350 3.500 ;
        RECT 44.680 3.330 44.850 3.500 ;
        RECT 48.880 5.830 49.050 6.000 ;
        RECT 49.380 5.830 49.550 6.000 ;
        RECT 49.880 5.830 50.050 6.000 ;
        RECT 50.380 5.830 50.550 6.000 ;
        RECT 50.880 5.830 51.050 6.000 ;
        RECT 51.380 5.830 51.550 6.000 ;
        RECT 48.880 5.330 49.050 5.500 ;
        RECT 49.380 5.330 49.550 5.500 ;
        RECT 49.880 5.330 50.050 5.500 ;
        RECT 50.380 5.330 50.550 5.500 ;
        RECT 50.880 5.330 51.050 5.500 ;
        RECT 51.380 5.330 51.550 5.500 ;
        RECT 48.880 4.830 49.050 5.000 ;
        RECT 49.380 4.830 49.550 5.000 ;
        RECT 49.880 4.830 50.050 5.000 ;
        RECT 50.380 4.830 50.550 5.000 ;
        RECT 50.880 4.830 51.050 5.000 ;
        RECT 51.380 4.830 51.550 5.000 ;
        RECT 48.880 4.330 49.050 4.500 ;
        RECT 49.380 4.330 49.550 4.500 ;
        RECT 49.880 4.330 50.050 4.500 ;
        RECT 50.380 4.330 50.550 4.500 ;
        RECT 50.880 4.330 51.050 4.500 ;
        RECT 51.380 4.330 51.550 4.500 ;
        RECT 48.880 3.830 49.050 4.000 ;
        RECT 49.380 3.830 49.550 4.000 ;
        RECT 49.880 3.830 50.050 4.000 ;
        RECT 50.380 3.830 50.550 4.000 ;
        RECT 50.880 3.830 51.050 4.000 ;
        RECT 51.380 3.830 51.550 4.000 ;
        RECT 48.880 3.330 49.050 3.500 ;
        RECT 49.380 3.330 49.550 3.500 ;
        RECT 49.880 3.330 50.050 3.500 ;
        RECT 50.380 3.330 50.550 3.500 ;
        RECT 50.880 3.330 51.050 3.500 ;
        RECT 51.380 3.330 51.550 3.500 ;
      LAYER met1 ;
        RECT 1.820 3.170 51.780 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 51.264000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 6.745 5.755 7.105 ;
        RECT 0.945 2.655 1.305 6.745 ;
        RECT 5.395 2.655 5.755 6.745 ;
        RECT 0.945 2.295 5.755 2.655 ;
        RECT 7.645 6.745 12.455 7.105 ;
        RECT 7.645 2.655 8.005 6.745 ;
        RECT 12.095 2.655 12.455 6.745 ;
        RECT 7.645 2.295 12.455 2.655 ;
        RECT 14.345 6.745 19.155 7.105 ;
        RECT 14.345 2.655 14.705 6.745 ;
        RECT 18.795 2.655 19.155 6.745 ;
        RECT 14.345 2.295 19.155 2.655 ;
        RECT 21.045 6.745 25.855 7.105 ;
        RECT 21.045 2.655 21.405 6.745 ;
        RECT 25.495 2.655 25.855 6.745 ;
        RECT 21.045 2.295 25.855 2.655 ;
        RECT 27.745 6.745 32.555 7.105 ;
        RECT 27.745 2.655 28.105 6.745 ;
        RECT 32.195 2.655 32.555 6.745 ;
        RECT 27.745 2.295 32.555 2.655 ;
        RECT 34.445 6.745 39.255 7.105 ;
        RECT 34.445 2.655 34.805 6.745 ;
        RECT 38.895 2.655 39.255 6.745 ;
        RECT 34.445 2.295 39.255 2.655 ;
        RECT 41.145 6.745 45.955 7.105 ;
        RECT 41.145 2.655 41.505 6.745 ;
        RECT 45.595 2.655 45.955 6.745 ;
        RECT 41.145 2.295 45.955 2.655 ;
        RECT 47.845 6.745 52.655 7.105 ;
        RECT 47.845 2.655 48.205 6.745 ;
        RECT 52.295 2.655 52.655 6.745 ;
        RECT 47.845 2.295 52.655 2.655 ;
      LAYER mcon ;
        RECT 1.050 6.850 1.220 7.020 ;
        RECT 1.500 6.850 1.670 7.020 ;
        RECT 1.950 6.850 2.120 7.020 ;
        RECT 2.400 6.850 2.570 7.020 ;
        RECT 2.850 6.850 3.020 7.020 ;
        RECT 3.300 6.850 3.470 7.020 ;
        RECT 3.750 6.850 3.920 7.020 ;
        RECT 4.200 6.850 4.370 7.020 ;
        RECT 4.650 6.850 4.820 7.020 ;
        RECT 5.100 6.850 5.270 7.020 ;
        RECT 5.550 6.850 5.720 7.020 ;
        RECT 7.750 6.850 7.920 7.020 ;
        RECT 8.200 6.850 8.370 7.020 ;
        RECT 8.650 6.850 8.820 7.020 ;
        RECT 9.100 6.850 9.270 7.020 ;
        RECT 9.550 6.850 9.720 7.020 ;
        RECT 10.000 6.850 10.170 7.020 ;
        RECT 10.450 6.850 10.620 7.020 ;
        RECT 10.900 6.850 11.070 7.020 ;
        RECT 11.350 6.850 11.520 7.020 ;
        RECT 11.800 6.850 11.970 7.020 ;
        RECT 12.250 6.850 12.420 7.020 ;
        RECT 14.450 6.850 14.620 7.020 ;
        RECT 14.900 6.850 15.070 7.020 ;
        RECT 15.350 6.850 15.520 7.020 ;
        RECT 15.800 6.850 15.970 7.020 ;
        RECT 16.250 6.850 16.420 7.020 ;
        RECT 16.700 6.850 16.870 7.020 ;
        RECT 17.150 6.850 17.320 7.020 ;
        RECT 17.600 6.850 17.770 7.020 ;
        RECT 18.050 6.850 18.220 7.020 ;
        RECT 18.500 6.850 18.670 7.020 ;
        RECT 18.950 6.850 19.120 7.020 ;
        RECT 21.150 6.850 21.320 7.020 ;
        RECT 21.600 6.850 21.770 7.020 ;
        RECT 22.050 6.850 22.220 7.020 ;
        RECT 22.500 6.850 22.670 7.020 ;
        RECT 22.950 6.850 23.120 7.020 ;
        RECT 23.400 6.850 23.570 7.020 ;
        RECT 23.850 6.850 24.020 7.020 ;
        RECT 24.300 6.850 24.470 7.020 ;
        RECT 24.750 6.850 24.920 7.020 ;
        RECT 25.200 6.850 25.370 7.020 ;
        RECT 25.650 6.850 25.820 7.020 ;
        RECT 27.850 6.850 28.020 7.020 ;
        RECT 28.300 6.850 28.470 7.020 ;
        RECT 28.750 6.850 28.920 7.020 ;
        RECT 29.200 6.850 29.370 7.020 ;
        RECT 29.650 6.850 29.820 7.020 ;
        RECT 30.100 6.850 30.270 7.020 ;
        RECT 30.550 6.850 30.720 7.020 ;
        RECT 31.000 6.850 31.170 7.020 ;
        RECT 31.450 6.850 31.620 7.020 ;
        RECT 31.900 6.850 32.070 7.020 ;
        RECT 32.350 6.850 32.520 7.020 ;
        RECT 34.550 6.850 34.720 7.020 ;
        RECT 35.000 6.850 35.170 7.020 ;
        RECT 35.450 6.850 35.620 7.020 ;
        RECT 35.900 6.850 36.070 7.020 ;
        RECT 36.350 6.850 36.520 7.020 ;
        RECT 36.800 6.850 36.970 7.020 ;
        RECT 37.250 6.850 37.420 7.020 ;
        RECT 37.700 6.850 37.870 7.020 ;
        RECT 38.150 6.850 38.320 7.020 ;
        RECT 38.600 6.850 38.770 7.020 ;
        RECT 39.050 6.850 39.220 7.020 ;
        RECT 41.250 6.850 41.420 7.020 ;
        RECT 41.700 6.850 41.870 7.020 ;
        RECT 42.150 6.850 42.320 7.020 ;
        RECT 42.600 6.850 42.770 7.020 ;
        RECT 43.050 6.850 43.220 7.020 ;
        RECT 43.500 6.850 43.670 7.020 ;
        RECT 43.950 6.850 44.120 7.020 ;
        RECT 44.400 6.850 44.570 7.020 ;
        RECT 44.850 6.850 45.020 7.020 ;
        RECT 45.300 6.850 45.470 7.020 ;
        RECT 45.750 6.850 45.920 7.020 ;
        RECT 47.950 6.850 48.120 7.020 ;
        RECT 48.400 6.850 48.570 7.020 ;
        RECT 48.850 6.850 49.020 7.020 ;
        RECT 49.300 6.850 49.470 7.020 ;
        RECT 49.750 6.850 49.920 7.020 ;
        RECT 50.200 6.850 50.370 7.020 ;
        RECT 50.650 6.850 50.820 7.020 ;
        RECT 51.100 6.850 51.270 7.020 ;
        RECT 51.550 6.850 51.720 7.020 ;
        RECT 52.000 6.850 52.170 7.020 ;
        RECT 52.450 6.850 52.620 7.020 ;
      LAYER met1 ;
        RECT 0.950 6.750 52.650 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 107.630394 ;
    PORT
      LAYER pwell ;
        RECT 0.000 7.285 53.600 8.050 ;
        RECT 0.000 2.115 0.765 7.285 ;
        RECT 5.935 2.115 7.465 7.285 ;
        RECT 12.635 2.115 14.165 7.285 ;
        RECT 19.335 2.115 20.865 7.285 ;
        RECT 26.035 2.115 27.565 7.285 ;
        RECT 32.735 2.115 34.265 7.285 ;
        RECT 39.435 2.115 40.965 7.285 ;
        RECT 46.135 2.115 47.665 7.285 ;
        RECT 52.835 2.115 53.600 7.285 ;
        RECT 0.000 1.350 53.600 2.115 ;
      LAYER li1 ;
        RECT 0.130 7.425 53.470 7.920 ;
        RECT 0.130 1.975 0.625 7.425 ;
        RECT 6.075 1.975 7.325 7.425 ;
        RECT 12.775 1.975 14.025 7.425 ;
        RECT 19.475 1.975 20.725 7.425 ;
        RECT 26.175 1.975 27.425 7.425 ;
        RECT 32.875 1.975 34.125 7.425 ;
        RECT 39.575 1.975 40.825 7.425 ;
        RECT 46.275 1.975 47.525 7.425 ;
        RECT 52.975 1.975 53.470 7.425 ;
        RECT 0.130 1.480 53.470 1.975 ;
      LAYER mcon ;
        RECT 0.230 7.650 0.400 7.820 ;
        RECT 0.680 7.650 0.850 7.820 ;
        RECT 1.130 7.650 1.300 7.820 ;
        RECT 1.580 7.650 1.750 7.820 ;
        RECT 2.030 7.650 2.200 7.820 ;
        RECT 2.480 7.650 2.650 7.820 ;
        RECT 2.930 7.650 3.100 7.820 ;
        RECT 3.380 7.650 3.550 7.820 ;
        RECT 3.830 7.650 4.000 7.820 ;
        RECT 4.280 7.650 4.450 7.820 ;
        RECT 4.730 7.650 4.900 7.820 ;
        RECT 5.180 7.650 5.350 7.820 ;
        RECT 5.630 7.650 5.800 7.820 ;
        RECT 6.080 7.650 6.250 7.820 ;
        RECT 6.930 7.650 7.100 7.820 ;
        RECT 7.380 7.650 7.550 7.820 ;
        RECT 7.830 7.650 8.000 7.820 ;
        RECT 8.280 7.650 8.450 7.820 ;
        RECT 8.730 7.650 8.900 7.820 ;
        RECT 9.180 7.650 9.350 7.820 ;
        RECT 9.630 7.650 9.800 7.820 ;
        RECT 10.080 7.650 10.250 7.820 ;
        RECT 10.530 7.650 10.700 7.820 ;
        RECT 10.980 7.650 11.150 7.820 ;
        RECT 11.430 7.650 11.600 7.820 ;
        RECT 11.880 7.650 12.050 7.820 ;
        RECT 12.330 7.650 12.500 7.820 ;
        RECT 12.780 7.650 12.950 7.820 ;
        RECT 13.630 7.650 13.800 7.820 ;
        RECT 14.080 7.650 14.250 7.820 ;
        RECT 14.530 7.650 14.700 7.820 ;
        RECT 14.980 7.650 15.150 7.820 ;
        RECT 15.430 7.650 15.600 7.820 ;
        RECT 15.880 7.650 16.050 7.820 ;
        RECT 16.330 7.650 16.500 7.820 ;
        RECT 16.780 7.650 16.950 7.820 ;
        RECT 17.230 7.650 17.400 7.820 ;
        RECT 17.680 7.650 17.850 7.820 ;
        RECT 18.130 7.650 18.300 7.820 ;
        RECT 18.580 7.650 18.750 7.820 ;
        RECT 19.030 7.650 19.200 7.820 ;
        RECT 19.480 7.650 19.650 7.820 ;
        RECT 20.330 7.650 20.500 7.820 ;
        RECT 20.780 7.650 20.950 7.820 ;
        RECT 21.230 7.650 21.400 7.820 ;
        RECT 21.680 7.650 21.850 7.820 ;
        RECT 22.130 7.650 22.300 7.820 ;
        RECT 22.580 7.650 22.750 7.820 ;
        RECT 23.030 7.650 23.200 7.820 ;
        RECT 23.480 7.650 23.650 7.820 ;
        RECT 23.930 7.650 24.100 7.820 ;
        RECT 24.380 7.650 24.550 7.820 ;
        RECT 24.830 7.650 25.000 7.820 ;
        RECT 25.280 7.650 25.450 7.820 ;
        RECT 25.730 7.650 25.900 7.820 ;
        RECT 26.180 7.650 26.350 7.820 ;
        RECT 27.030 7.650 27.200 7.820 ;
        RECT 27.480 7.650 27.650 7.820 ;
        RECT 27.930 7.650 28.100 7.820 ;
        RECT 28.380 7.650 28.550 7.820 ;
        RECT 28.830 7.650 29.000 7.820 ;
        RECT 29.280 7.650 29.450 7.820 ;
        RECT 29.730 7.650 29.900 7.820 ;
        RECT 30.180 7.650 30.350 7.820 ;
        RECT 30.630 7.650 30.800 7.820 ;
        RECT 31.080 7.650 31.250 7.820 ;
        RECT 31.530 7.650 31.700 7.820 ;
        RECT 31.980 7.650 32.150 7.820 ;
        RECT 32.430 7.650 32.600 7.820 ;
        RECT 32.880 7.650 33.050 7.820 ;
        RECT 33.730 7.650 33.900 7.820 ;
        RECT 34.180 7.650 34.350 7.820 ;
        RECT 34.630 7.650 34.800 7.820 ;
        RECT 35.080 7.650 35.250 7.820 ;
        RECT 35.530 7.650 35.700 7.820 ;
        RECT 35.980 7.650 36.150 7.820 ;
        RECT 36.430 7.650 36.600 7.820 ;
        RECT 36.880 7.650 37.050 7.820 ;
        RECT 37.330 7.650 37.500 7.820 ;
        RECT 37.780 7.650 37.950 7.820 ;
        RECT 38.230 7.650 38.400 7.820 ;
        RECT 38.680 7.650 38.850 7.820 ;
        RECT 39.130 7.650 39.300 7.820 ;
        RECT 39.580 7.650 39.750 7.820 ;
        RECT 40.430 7.650 40.600 7.820 ;
        RECT 40.880 7.650 41.050 7.820 ;
        RECT 41.330 7.650 41.500 7.820 ;
        RECT 41.780 7.650 41.950 7.820 ;
        RECT 42.230 7.650 42.400 7.820 ;
        RECT 42.680 7.650 42.850 7.820 ;
        RECT 43.130 7.650 43.300 7.820 ;
        RECT 43.580 7.650 43.750 7.820 ;
        RECT 44.030 7.650 44.200 7.820 ;
        RECT 44.480 7.650 44.650 7.820 ;
        RECT 44.930 7.650 45.100 7.820 ;
        RECT 45.380 7.650 45.550 7.820 ;
        RECT 45.830 7.650 46.000 7.820 ;
        RECT 46.280 7.650 46.450 7.820 ;
        RECT 47.130 7.650 47.300 7.820 ;
        RECT 47.580 7.650 47.750 7.820 ;
        RECT 48.030 7.650 48.200 7.820 ;
        RECT 48.480 7.650 48.650 7.820 ;
        RECT 48.930 7.650 49.100 7.820 ;
        RECT 49.380 7.650 49.550 7.820 ;
        RECT 49.830 7.650 50.000 7.820 ;
        RECT 50.280 7.650 50.450 7.820 ;
        RECT 50.730 7.650 50.900 7.820 ;
        RECT 51.180 7.650 51.350 7.820 ;
        RECT 51.630 7.650 51.800 7.820 ;
        RECT 52.080 7.650 52.250 7.820 ;
        RECT 52.530 7.650 52.700 7.820 ;
        RECT 52.980 7.650 53.150 7.820 ;
      LAYER met1 ;
        RECT 0.130 7.500 53.470 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 53.600 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 1.850 9.250 2.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 3.850 9.250 4.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 5.850 9.250 6.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 7.850 9.250 8.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 9.850 9.250 10.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 11.850 9.250 12.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 13.850 9.250 14.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 15.850 9.250 16.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 17.850 9.250 18.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
        RECT 19.850 9.250 20.150 9.550 ;
        RECT 20.850 9.250 21.150 9.550 ;
        RECT 21.850 9.250 22.150 9.550 ;
        RECT 22.850 9.250 23.150 9.550 ;
        RECT 23.850 9.250 24.150 9.550 ;
        RECT 24.850 9.250 25.150 9.550 ;
        RECT 25.850 9.250 26.150 9.550 ;
        RECT 26.850 9.250 27.150 9.550 ;
        RECT 27.850 9.250 28.150 9.550 ;
        RECT 28.850 9.250 29.150 9.550 ;
        RECT 29.850 9.250 30.150 9.550 ;
        RECT 30.850 9.250 31.150 9.550 ;
        RECT 31.850 9.250 32.150 9.550 ;
        RECT 32.850 9.250 33.150 9.550 ;
        RECT 33.850 9.250 34.150 9.550 ;
        RECT 34.850 9.250 35.150 9.550 ;
        RECT 35.850 9.250 36.150 9.550 ;
        RECT 36.850 9.250 37.150 9.550 ;
        RECT 37.850 9.250 38.150 9.550 ;
        RECT 38.850 9.250 39.150 9.550 ;
        RECT 39.850 9.250 40.150 9.550 ;
        RECT 40.850 9.250 41.150 9.550 ;
        RECT 41.850 9.250 42.150 9.550 ;
        RECT 42.850 9.250 43.150 9.550 ;
        RECT 43.850 9.250 44.150 9.550 ;
        RECT 44.850 9.250 45.150 9.550 ;
        RECT 45.850 9.250 46.150 9.550 ;
        RECT 46.850 9.250 47.150 9.550 ;
        RECT 47.850 9.250 48.150 9.550 ;
        RECT 48.850 9.250 49.150 9.550 ;
        RECT 49.850 9.250 50.150 9.550 ;
        RECT 50.850 9.250 51.150 9.550 ;
        RECT 51.850 9.250 52.150 9.550 ;
        RECT 52.850 9.250 53.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 53.600 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 53.600 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.850 -0.150 21.150 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.850 -0.150 23.150 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.850 -0.150 25.150 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.850 -0.150 27.150 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.850 -0.150 29.150 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.850 -0.150 31.150 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.850 -0.150 33.150 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.850 -0.150 35.150 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.850 -0.150 37.150 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.850 -0.150 39.150 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.850 -0.150 41.150 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.850 -0.150 43.150 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.850 -0.150 45.150 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
        RECT 46.850 -0.150 47.150 0.150 ;
        RECT 47.850 -0.150 48.150 0.150 ;
        RECT 48.850 -0.150 49.150 0.150 ;
        RECT 49.850 -0.150 50.150 0.150 ;
        RECT 50.850 -0.150 51.150 0.150 ;
        RECT 51.850 -0.150 52.150 0.150 ;
        RECT 52.850 -0.150 53.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 53.600 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_8
END LIBRARY

