magic
tech sky130A
magscale 1 2
timestamp 1658609782
<< nwell >>
rect 130 1707 5756 1940
rect 130 1000 5757 1707
rect 131 293 5757 1000
<< pmoslvt >>
rect 225 355 625 1645
rect 683 355 1083 1645
rect 1141 355 1541 1645
rect 1599 355 1999 1645
rect 2057 355 2457 1645
rect 2515 355 2915 1645
rect 2973 355 3373 1645
rect 3431 355 3831 1645
rect 3889 355 4289 1645
rect 4347 355 4747 1645
rect 4805 355 5205 1645
rect 5263 355 5663 1645
<< pdiff >>
rect 167 1633 225 1645
rect 167 367 179 1633
rect 213 367 225 1633
rect 167 355 225 367
rect 625 1633 683 1645
rect 625 367 637 1633
rect 671 367 683 1633
rect 625 355 683 367
rect 1083 1633 1141 1645
rect 1083 367 1095 1633
rect 1129 367 1141 1633
rect 1083 355 1141 367
rect 1541 1633 1599 1645
rect 1541 367 1553 1633
rect 1587 367 1599 1633
rect 1541 355 1599 367
rect 1999 1633 2057 1645
rect 1999 367 2011 1633
rect 2045 367 2057 1633
rect 1999 355 2057 367
rect 2457 1633 2515 1645
rect 2457 367 2469 1633
rect 2503 367 2515 1633
rect 2457 355 2515 367
rect 2915 1633 2973 1645
rect 2915 367 2927 1633
rect 2961 367 2973 1633
rect 2915 355 2973 367
rect 3373 1633 3431 1645
rect 3373 367 3385 1633
rect 3419 367 3431 1633
rect 3373 355 3431 367
rect 3831 1633 3889 1645
rect 3831 367 3843 1633
rect 3877 367 3889 1633
rect 3831 355 3889 367
rect 4289 1633 4347 1645
rect 4289 367 4301 1633
rect 4335 367 4347 1633
rect 4289 355 4347 367
rect 4747 1633 4805 1645
rect 4747 367 4759 1633
rect 4793 367 4805 1633
rect 4747 355 4805 367
rect 5205 1633 5263 1645
rect 5205 367 5217 1633
rect 5251 367 5263 1633
rect 5205 355 5263 367
rect 5663 1633 5721 1645
rect 5663 367 5675 1633
rect 5709 367 5721 1633
rect 5663 355 5721 367
<< pdiffc >>
rect 179 367 213 1633
rect 637 367 671 1633
rect 1095 367 1129 1633
rect 1553 367 1587 1633
rect 2011 367 2045 1633
rect 2469 367 2503 1633
rect 2927 367 2961 1633
rect 3385 367 3419 1633
rect 3843 367 3877 1633
rect 4301 367 4335 1633
rect 4759 367 4793 1633
rect 5217 367 5251 1633
rect 5675 367 5709 1633
<< poly >>
rect 225 1645 625 1671
rect 683 1645 1083 1671
rect 1141 1645 1541 1671
rect 1599 1645 1999 1671
rect 2057 1645 2457 1671
rect 2515 1645 2915 1671
rect 2973 1645 3373 1671
rect 3431 1645 3831 1671
rect 3889 1645 4289 1671
rect 4347 1645 4747 1671
rect 4805 1645 5205 1671
rect 5263 1645 5663 1671
rect 225 329 625 355
rect 683 329 1083 355
rect 1141 329 1541 355
rect 1599 329 1999 355
rect 2057 329 2457 355
rect 2515 329 2915 355
rect 2973 329 3373 355
rect 3431 329 3831 355
rect 3889 329 4289 355
rect 4347 329 4747 355
rect 4805 329 5205 355
rect 5263 329 5663 355
rect 370 182 490 329
rect 826 182 946 329
rect 1282 182 1402 329
rect 1738 182 1858 329
rect 2194 182 2314 329
rect 2650 182 2770 329
rect 3106 182 3226 329
rect 3562 182 3682 329
rect 4018 182 4138 329
rect 4474 182 4594 329
rect 4930 182 5050 329
rect 5386 182 5506 329
rect 130 162 5756 182
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3100 162
rect 3160 102 3500 162
rect 3560 102 3900 162
rect 3960 102 4300 162
rect 4360 102 4700 162
rect 4760 102 5100 162
rect 5160 102 5500 162
rect 5560 102 5756 162
rect 130 82 5756 102
<< polycont >>
rect 300 102 360 162
rect 700 102 760 162
rect 1100 102 1160 162
rect 1500 102 1560 162
rect 1900 102 1960 162
rect 2300 102 2360 162
rect 2700 102 2760 162
rect 3100 102 3160 162
rect 3500 102 3560 162
rect 3900 102 3960 162
rect 4300 102 4360 162
rect 4700 102 4760 162
rect 5100 102 5160 162
rect 5500 102 5560 162
<< locali >>
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3100 1910
rect 3160 1850 3500 1910
rect 3560 1850 3900 1910
rect 3960 1850 4300 1910
rect 4360 1850 4700 1910
rect 4760 1850 5100 1910
rect 5160 1850 5500 1910
rect 5560 1850 5756 1910
rect 130 1730 5756 1790
rect 635 1649 669 1730
rect 1551 1649 1585 1730
rect 2467 1649 2501 1730
rect 3383 1649 3417 1730
rect 4299 1649 4333 1730
rect 5215 1649 5249 1730
rect 179 1633 213 1649
rect 177 367 179 372
rect 635 1633 671 1649
rect 635 1626 637 1633
rect 177 351 213 367
rect 1095 1633 1129 1649
rect 637 351 671 367
rect 1093 367 1095 372
rect 1551 1633 1587 1649
rect 1551 1626 1553 1633
rect 1093 351 1129 367
rect 2011 1633 2045 1649
rect 1553 351 1587 367
rect 2009 367 2011 372
rect 2467 1633 2503 1649
rect 2467 1626 2469 1633
rect 2009 351 2045 367
rect 2927 1633 2961 1649
rect 2469 351 2503 367
rect 2925 367 2927 372
rect 3383 1633 3419 1649
rect 3383 1626 3385 1633
rect 2925 351 2961 367
rect 3843 1633 3877 1649
rect 3385 351 3419 367
rect 3841 367 3843 372
rect 4299 1633 4335 1649
rect 4299 1626 4301 1633
rect 3841 351 3877 367
rect 4759 1633 4793 1649
rect 4301 351 4335 367
rect 4757 367 4759 372
rect 5215 1633 5251 1649
rect 5215 1626 5217 1633
rect 4757 351 4793 367
rect 5675 1633 5709 1649
rect 5217 351 5251 367
rect 5673 367 5675 372
rect 5673 351 5709 367
rect 177 270 211 351
rect 1093 270 1127 351
rect 2009 270 2043 351
rect 2925 270 2959 351
rect 3841 270 3875 351
rect 4757 270 4791 351
rect 5673 270 5707 351
rect 130 210 5756 270
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3100 162
rect 3160 102 3500 162
rect 3560 102 3900 162
rect 3960 102 4300 162
rect 4360 102 4700 162
rect 4760 102 5100 162
rect 5160 102 5500 162
rect 5560 102 5756 162
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3100 30
rect 3160 -30 3500 30
rect 3560 -30 3900 30
rect 3960 -30 4300 30
rect 4360 -30 4700 30
rect 4760 -30 5100 30
rect 5160 -30 5500 30
rect 5560 -30 5756 30
<< viali >>
rect 300 1850 360 1910
rect 700 1850 760 1910
rect 1100 1850 1160 1910
rect 1500 1850 1560 1910
rect 1900 1850 1960 1910
rect 2300 1850 2360 1910
rect 2700 1850 2760 1910
rect 3100 1850 3160 1910
rect 3500 1850 3560 1910
rect 3900 1850 3960 1910
rect 4300 1850 4360 1910
rect 4700 1850 4760 1910
rect 5100 1850 5160 1910
rect 5500 1850 5560 1910
rect 179 367 213 1633
rect 637 367 671 1633
rect 1095 367 1129 1633
rect 1553 367 1587 1633
rect 2011 367 2045 1633
rect 2469 367 2503 1633
rect 2927 367 2961 1633
rect 3385 367 3419 1633
rect 3843 367 3877 1633
rect 4301 367 4335 1633
rect 4759 367 4793 1633
rect 5217 367 5251 1633
rect 5675 367 5709 1633
rect 300 -30 360 30
rect 700 -30 760 30
rect 1100 -30 1160 30
rect 1500 -30 1560 30
rect 1900 -30 1960 30
rect 2300 -30 2360 30
rect 2700 -30 2760 30
rect 3100 -30 3160 30
rect 3500 -30 3560 30
rect 3900 -30 3960 30
rect 4300 -30 4360 30
rect 4700 -30 4760 30
rect 5100 -30 5160 30
rect 5500 -30 5560 30
<< metal1 >>
rect 130 1910 5756 1940
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3100 1910
rect 3160 1850 3500 1910
rect 3560 1850 3900 1910
rect 3960 1850 4300 1910
rect 4360 1850 4700 1910
rect 4760 1850 5100 1910
rect 5160 1850 5500 1910
rect 5560 1850 5756 1910
rect 130 1820 5756 1850
rect 173 1633 219 1645
rect 173 367 179 1633
rect 213 367 219 1633
rect 173 355 219 367
rect 631 1633 677 1645
rect 631 367 637 1633
rect 671 367 677 1633
rect 631 355 677 367
rect 1089 1633 1135 1645
rect 1089 367 1095 1633
rect 1129 367 1135 1633
rect 1089 355 1135 367
rect 1547 1633 1593 1645
rect 1547 367 1553 1633
rect 1587 367 1593 1633
rect 1547 355 1593 367
rect 2005 1633 2051 1645
rect 2005 367 2011 1633
rect 2045 367 2051 1633
rect 2005 355 2051 367
rect 2463 1633 2509 1645
rect 2463 367 2469 1633
rect 2503 367 2509 1633
rect 2463 355 2509 367
rect 2921 1633 2967 1645
rect 2921 367 2927 1633
rect 2961 367 2967 1633
rect 2921 355 2967 367
rect 3379 1633 3425 1645
rect 3379 367 3385 1633
rect 3419 367 3425 1633
rect 3379 355 3425 367
rect 3837 1633 3883 1645
rect 3837 367 3843 1633
rect 3877 367 3883 1633
rect 3837 355 3883 367
rect 4295 1633 4341 1645
rect 4295 367 4301 1633
rect 4335 367 4341 1633
rect 4295 355 4341 367
rect 4753 1633 4799 1645
rect 4753 367 4759 1633
rect 4793 367 4799 1633
rect 4753 355 4799 367
rect 5211 1633 5257 1645
rect 5211 367 5217 1633
rect 5251 367 5257 1633
rect 5211 355 5257 367
rect 5669 1633 5715 1645
rect 5669 367 5675 1633
rect 5709 367 5715 1633
rect 5669 355 5715 367
rect 130 30 5756 60
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3100 30
rect 3160 -30 3500 30
rect 3560 -30 3900 30
rect 3960 -30 4300 30
rect 4360 -30 4700 30
rect 4760 -30 5100 30
rect 5160 -30 5500 30
rect 5560 -30 5756 30
rect 130 -60 5756 -30
<< labels >>
flabel metal1 130 1850 190 1910 1 FreeSans 480 0 0 0 VPWR
port 4 n power bidirectional
flabel space 120 1850 180 1910 1 FreeSans 480 0 0 0 VPB
flabel metal1 130 -30 190 30 1 FreeSans 480 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 5696 1730 5756 1790 1 FreeSans 480 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 5696 210 5756 270 1 FreeSans 480 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 5696 102 5756 162 1 FreeSans 480 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5963 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
